module sincos (
	icos,  //out
	qsin,  //out
	t,	   //in
	i,
	q
);

output [8:0] icos;
output [8:0] qsin;

input [4:0] t;
input [`IQMSB:0] i;
input [`IQMSB:0] q;

reg signed [8:0] icos_lut [0:8191];
reg signed [8:0] qsin_lut [0:8191];

// address [12:5] is the multiplier:
//	 0:-1, (127,128)=~0, 255=1
// address [4:0] is t

assign icos=icos_lut[{i,t}];
assign qsin=qsin_lut[{q,t}];

// generated with iq_lut.pl
initial begin
	qsin_lut[0000] =  9'sd0;
	icos_lut[0000] = -9'sd255;
	qsin_lut[0001] = -9'sd50;
	icos_lut[0001] = -9'sd250;
	qsin_lut[0002] = -9'sd98;
	icos_lut[0002] = -9'sd236;
	qsin_lut[0003] = -9'sd142;
	icos_lut[0003] = -9'sd212;
	qsin_lut[0004] = -9'sd180;
	icos_lut[0004] = -9'sd180;
	qsin_lut[0005] = -9'sd212;
	icos_lut[0005] = -9'sd142;
	qsin_lut[0006] = -9'sd236;
	icos_lut[0006] = -9'sd98;
	qsin_lut[0007] = -9'sd250;
	icos_lut[0007] = -9'sd50;
	qsin_lut[0008] = -9'sd255;
	icos_lut[0008] = -9'sd0;
	qsin_lut[0009] = -9'sd250;
	icos_lut[0009] =  9'sd50;
	qsin_lut[0010] = -9'sd236;
	icos_lut[0010] =  9'sd98;
	qsin_lut[0011] = -9'sd212;
	icos_lut[0011] =  9'sd142;
	qsin_lut[0012] = -9'sd180;
	icos_lut[0012] =  9'sd180;
	qsin_lut[0013] = -9'sd142;
	icos_lut[0013] =  9'sd212;
	qsin_lut[0014] = -9'sd98;
	icos_lut[0014] =  9'sd236;
	qsin_lut[0015] = -9'sd50;
	icos_lut[0015] =  9'sd250;
	qsin_lut[0016] = -9'sd0;
	icos_lut[0016] =  9'sd255;
	qsin_lut[0017] =  9'sd50;
	icos_lut[0017] =  9'sd250;
	qsin_lut[0018] =  9'sd98;
	icos_lut[0018] =  9'sd236;
	qsin_lut[0019] =  9'sd142;
	icos_lut[0019] =  9'sd212;
	qsin_lut[0020] =  9'sd180;
	icos_lut[0020] =  9'sd180;
	qsin_lut[0021] =  9'sd212;
	icos_lut[0021] =  9'sd142;
	qsin_lut[0022] =  9'sd236;
	icos_lut[0022] =  9'sd98;
	qsin_lut[0023] =  9'sd250;
	icos_lut[0023] =  9'sd50;
	qsin_lut[0024] =  9'sd255;
	icos_lut[0024] =  9'sd0;
	qsin_lut[0025] =  9'sd250;
	icos_lut[0025] = -9'sd50;
	qsin_lut[0026] =  9'sd236;
	icos_lut[0026] = -9'sd98;
	qsin_lut[0027] =  9'sd212;
	icos_lut[0027] = -9'sd142;
	qsin_lut[0028] =  9'sd180;
	icos_lut[0028] = -9'sd180;
	qsin_lut[0029] =  9'sd142;
	icos_lut[0029] = -9'sd212;
	qsin_lut[0030] =  9'sd98;
	icos_lut[0030] = -9'sd236;
	qsin_lut[0031] =  9'sd50;
	icos_lut[0031] = -9'sd250;
	qsin_lut[0032] =  9'sd0;
	icos_lut[0032] = -9'sd253;
	qsin_lut[0033] = -9'sd49;
	icos_lut[0033] = -9'sd248;
	qsin_lut[0034] = -9'sd97;
	icos_lut[0034] = -9'sd234;
	qsin_lut[0035] = -9'sd141;
	icos_lut[0035] = -9'sd210;
	qsin_lut[0036] = -9'sd179;
	icos_lut[0036] = -9'sd179;
	qsin_lut[0037] = -9'sd210;
	icos_lut[0037] = -9'sd141;
	qsin_lut[0038] = -9'sd234;
	icos_lut[0038] = -9'sd97;
	qsin_lut[0039] = -9'sd248;
	icos_lut[0039] = -9'sd49;
	qsin_lut[0040] = -9'sd253;
	icos_lut[0040] = -9'sd0;
	qsin_lut[0041] = -9'sd248;
	icos_lut[0041] =  9'sd49;
	qsin_lut[0042] = -9'sd234;
	icos_lut[0042] =  9'sd97;
	qsin_lut[0043] = -9'sd210;
	icos_lut[0043] =  9'sd141;
	qsin_lut[0044] = -9'sd179;
	icos_lut[0044] =  9'sd179;
	qsin_lut[0045] = -9'sd141;
	icos_lut[0045] =  9'sd210;
	qsin_lut[0046] = -9'sd97;
	icos_lut[0046] =  9'sd234;
	qsin_lut[0047] = -9'sd49;
	icos_lut[0047] =  9'sd248;
	qsin_lut[0048] = -9'sd0;
	icos_lut[0048] =  9'sd253;
	qsin_lut[0049] =  9'sd49;
	icos_lut[0049] =  9'sd248;
	qsin_lut[0050] =  9'sd97;
	icos_lut[0050] =  9'sd234;
	qsin_lut[0051] =  9'sd141;
	icos_lut[0051] =  9'sd210;
	qsin_lut[0052] =  9'sd179;
	icos_lut[0052] =  9'sd179;
	qsin_lut[0053] =  9'sd210;
	icos_lut[0053] =  9'sd141;
	qsin_lut[0054] =  9'sd234;
	icos_lut[0054] =  9'sd97;
	qsin_lut[0055] =  9'sd248;
	icos_lut[0055] =  9'sd49;
	qsin_lut[0056] =  9'sd253;
	icos_lut[0056] =  9'sd0;
	qsin_lut[0057] =  9'sd248;
	icos_lut[0057] = -9'sd49;
	qsin_lut[0058] =  9'sd234;
	icos_lut[0058] = -9'sd97;
	qsin_lut[0059] =  9'sd210;
	icos_lut[0059] = -9'sd141;
	qsin_lut[0060] =  9'sd179;
	icos_lut[0060] = -9'sd179;
	qsin_lut[0061] =  9'sd141;
	icos_lut[0061] = -9'sd210;
	qsin_lut[0062] =  9'sd97;
	icos_lut[0062] = -9'sd234;
	qsin_lut[0063] =  9'sd49;
	icos_lut[0063] = -9'sd248;
	qsin_lut[0064] =  9'sd0;
	icos_lut[0064] = -9'sd251;
	qsin_lut[0065] = -9'sd49;
	icos_lut[0065] = -9'sd246;
	qsin_lut[0066] = -9'sd96;
	icos_lut[0066] = -9'sd232;
	qsin_lut[0067] = -9'sd139;
	icos_lut[0067] = -9'sd209;
	qsin_lut[0068] = -9'sd177;
	icos_lut[0068] = -9'sd177;
	qsin_lut[0069] = -9'sd209;
	icos_lut[0069] = -9'sd139;
	qsin_lut[0070] = -9'sd232;
	icos_lut[0070] = -9'sd96;
	qsin_lut[0071] = -9'sd246;
	icos_lut[0071] = -9'sd49;
	qsin_lut[0072] = -9'sd251;
	icos_lut[0072] = -9'sd0;
	qsin_lut[0073] = -9'sd246;
	icos_lut[0073] =  9'sd49;
	qsin_lut[0074] = -9'sd232;
	icos_lut[0074] =  9'sd96;
	qsin_lut[0075] = -9'sd209;
	icos_lut[0075] =  9'sd139;
	qsin_lut[0076] = -9'sd177;
	icos_lut[0076] =  9'sd177;
	qsin_lut[0077] = -9'sd139;
	icos_lut[0077] =  9'sd209;
	qsin_lut[0078] = -9'sd96;
	icos_lut[0078] =  9'sd232;
	qsin_lut[0079] = -9'sd49;
	icos_lut[0079] =  9'sd246;
	qsin_lut[0080] = -9'sd0;
	icos_lut[0080] =  9'sd251;
	qsin_lut[0081] =  9'sd49;
	icos_lut[0081] =  9'sd246;
	qsin_lut[0082] =  9'sd96;
	icos_lut[0082] =  9'sd232;
	qsin_lut[0083] =  9'sd139;
	icos_lut[0083] =  9'sd209;
	qsin_lut[0084] =  9'sd177;
	icos_lut[0084] =  9'sd177;
	qsin_lut[0085] =  9'sd209;
	icos_lut[0085] =  9'sd139;
	qsin_lut[0086] =  9'sd232;
	icos_lut[0086] =  9'sd96;
	qsin_lut[0087] =  9'sd246;
	icos_lut[0087] =  9'sd49;
	qsin_lut[0088] =  9'sd251;
	icos_lut[0088] =  9'sd0;
	qsin_lut[0089] =  9'sd246;
	icos_lut[0089] = -9'sd49;
	qsin_lut[0090] =  9'sd232;
	icos_lut[0090] = -9'sd96;
	qsin_lut[0091] =  9'sd209;
	icos_lut[0091] = -9'sd139;
	qsin_lut[0092] =  9'sd177;
	icos_lut[0092] = -9'sd177;
	qsin_lut[0093] =  9'sd139;
	icos_lut[0093] = -9'sd209;
	qsin_lut[0094] =  9'sd96;
	icos_lut[0094] = -9'sd232;
	qsin_lut[0095] =  9'sd49;
	icos_lut[0095] = -9'sd246;
	qsin_lut[0096] =  9'sd0;
	icos_lut[0096] = -9'sd249;
	qsin_lut[0097] = -9'sd49;
	icos_lut[0097] = -9'sd244;
	qsin_lut[0098] = -9'sd95;
	icos_lut[0098] = -9'sd230;
	qsin_lut[0099] = -9'sd138;
	icos_lut[0099] = -9'sd207;
	qsin_lut[0100] = -9'sd176;
	icos_lut[0100] = -9'sd176;
	qsin_lut[0101] = -9'sd207;
	icos_lut[0101] = -9'sd138;
	qsin_lut[0102] = -9'sd230;
	icos_lut[0102] = -9'sd95;
	qsin_lut[0103] = -9'sd244;
	icos_lut[0103] = -9'sd49;
	qsin_lut[0104] = -9'sd249;
	icos_lut[0104] = -9'sd0;
	qsin_lut[0105] = -9'sd244;
	icos_lut[0105] =  9'sd49;
	qsin_lut[0106] = -9'sd230;
	icos_lut[0106] =  9'sd95;
	qsin_lut[0107] = -9'sd207;
	icos_lut[0107] =  9'sd138;
	qsin_lut[0108] = -9'sd176;
	icos_lut[0108] =  9'sd176;
	qsin_lut[0109] = -9'sd138;
	icos_lut[0109] =  9'sd207;
	qsin_lut[0110] = -9'sd95;
	icos_lut[0110] =  9'sd230;
	qsin_lut[0111] = -9'sd49;
	icos_lut[0111] =  9'sd244;
	qsin_lut[0112] = -9'sd0;
	icos_lut[0112] =  9'sd249;
	qsin_lut[0113] =  9'sd49;
	icos_lut[0113] =  9'sd244;
	qsin_lut[0114] =  9'sd95;
	icos_lut[0114] =  9'sd230;
	qsin_lut[0115] =  9'sd138;
	icos_lut[0115] =  9'sd207;
	qsin_lut[0116] =  9'sd176;
	icos_lut[0116] =  9'sd176;
	qsin_lut[0117] =  9'sd207;
	icos_lut[0117] =  9'sd138;
	qsin_lut[0118] =  9'sd230;
	icos_lut[0118] =  9'sd95;
	qsin_lut[0119] =  9'sd244;
	icos_lut[0119] =  9'sd49;
	qsin_lut[0120] =  9'sd249;
	icos_lut[0120] =  9'sd0;
	qsin_lut[0121] =  9'sd244;
	icos_lut[0121] = -9'sd49;
	qsin_lut[0122] =  9'sd230;
	icos_lut[0122] = -9'sd95;
	qsin_lut[0123] =  9'sd207;
	icos_lut[0123] = -9'sd138;
	qsin_lut[0124] =  9'sd176;
	icos_lut[0124] = -9'sd176;
	qsin_lut[0125] =  9'sd138;
	icos_lut[0125] = -9'sd207;
	qsin_lut[0126] =  9'sd95;
	icos_lut[0126] = -9'sd230;
	qsin_lut[0127] =  9'sd49;
	icos_lut[0127] = -9'sd244;
	qsin_lut[0128] =  9'sd0;
	icos_lut[0128] = -9'sd247;
	qsin_lut[0129] = -9'sd48;
	icos_lut[0129] = -9'sd242;
	qsin_lut[0130] = -9'sd95;
	icos_lut[0130] = -9'sd228;
	qsin_lut[0131] = -9'sd137;
	icos_lut[0131] = -9'sd205;
	qsin_lut[0132] = -9'sd175;
	icos_lut[0132] = -9'sd175;
	qsin_lut[0133] = -9'sd205;
	icos_lut[0133] = -9'sd137;
	qsin_lut[0134] = -9'sd228;
	icos_lut[0134] = -9'sd95;
	qsin_lut[0135] = -9'sd242;
	icos_lut[0135] = -9'sd48;
	qsin_lut[0136] = -9'sd247;
	icos_lut[0136] = -9'sd0;
	qsin_lut[0137] = -9'sd242;
	icos_lut[0137] =  9'sd48;
	qsin_lut[0138] = -9'sd228;
	icos_lut[0138] =  9'sd95;
	qsin_lut[0139] = -9'sd205;
	icos_lut[0139] =  9'sd137;
	qsin_lut[0140] = -9'sd175;
	icos_lut[0140] =  9'sd175;
	qsin_lut[0141] = -9'sd137;
	icos_lut[0141] =  9'sd205;
	qsin_lut[0142] = -9'sd95;
	icos_lut[0142] =  9'sd228;
	qsin_lut[0143] = -9'sd48;
	icos_lut[0143] =  9'sd242;
	qsin_lut[0144] = -9'sd0;
	icos_lut[0144] =  9'sd247;
	qsin_lut[0145] =  9'sd48;
	icos_lut[0145] =  9'sd242;
	qsin_lut[0146] =  9'sd95;
	icos_lut[0146] =  9'sd228;
	qsin_lut[0147] =  9'sd137;
	icos_lut[0147] =  9'sd205;
	qsin_lut[0148] =  9'sd175;
	icos_lut[0148] =  9'sd175;
	qsin_lut[0149] =  9'sd205;
	icos_lut[0149] =  9'sd137;
	qsin_lut[0150] =  9'sd228;
	icos_lut[0150] =  9'sd95;
	qsin_lut[0151] =  9'sd242;
	icos_lut[0151] =  9'sd48;
	qsin_lut[0152] =  9'sd247;
	icos_lut[0152] =  9'sd0;
	qsin_lut[0153] =  9'sd242;
	icos_lut[0153] = -9'sd48;
	qsin_lut[0154] =  9'sd228;
	icos_lut[0154] = -9'sd95;
	qsin_lut[0155] =  9'sd205;
	icos_lut[0155] = -9'sd137;
	qsin_lut[0156] =  9'sd175;
	icos_lut[0156] = -9'sd175;
	qsin_lut[0157] =  9'sd137;
	icos_lut[0157] = -9'sd205;
	qsin_lut[0158] =  9'sd95;
	icos_lut[0158] = -9'sd228;
	qsin_lut[0159] =  9'sd48;
	icos_lut[0159] = -9'sd242;
	qsin_lut[0160] =  9'sd0;
	icos_lut[0160] = -9'sd245;
	qsin_lut[0161] = -9'sd48;
	icos_lut[0161] = -9'sd240;
	qsin_lut[0162] = -9'sd94;
	icos_lut[0162] = -9'sd226;
	qsin_lut[0163] = -9'sd136;
	icos_lut[0163] = -9'sd204;
	qsin_lut[0164] = -9'sd173;
	icos_lut[0164] = -9'sd173;
	qsin_lut[0165] = -9'sd204;
	icos_lut[0165] = -9'sd136;
	qsin_lut[0166] = -9'sd226;
	icos_lut[0166] = -9'sd94;
	qsin_lut[0167] = -9'sd240;
	icos_lut[0167] = -9'sd48;
	qsin_lut[0168] = -9'sd245;
	icos_lut[0168] = -9'sd0;
	qsin_lut[0169] = -9'sd240;
	icos_lut[0169] =  9'sd48;
	qsin_lut[0170] = -9'sd226;
	icos_lut[0170] =  9'sd94;
	qsin_lut[0171] = -9'sd204;
	icos_lut[0171] =  9'sd136;
	qsin_lut[0172] = -9'sd173;
	icos_lut[0172] =  9'sd173;
	qsin_lut[0173] = -9'sd136;
	icos_lut[0173] =  9'sd204;
	qsin_lut[0174] = -9'sd94;
	icos_lut[0174] =  9'sd226;
	qsin_lut[0175] = -9'sd48;
	icos_lut[0175] =  9'sd240;
	qsin_lut[0176] = -9'sd0;
	icos_lut[0176] =  9'sd245;
	qsin_lut[0177] =  9'sd48;
	icos_lut[0177] =  9'sd240;
	qsin_lut[0178] =  9'sd94;
	icos_lut[0178] =  9'sd226;
	qsin_lut[0179] =  9'sd136;
	icos_lut[0179] =  9'sd204;
	qsin_lut[0180] =  9'sd173;
	icos_lut[0180] =  9'sd173;
	qsin_lut[0181] =  9'sd204;
	icos_lut[0181] =  9'sd136;
	qsin_lut[0182] =  9'sd226;
	icos_lut[0182] =  9'sd94;
	qsin_lut[0183] =  9'sd240;
	icos_lut[0183] =  9'sd48;
	qsin_lut[0184] =  9'sd245;
	icos_lut[0184] =  9'sd0;
	qsin_lut[0185] =  9'sd240;
	icos_lut[0185] = -9'sd48;
	qsin_lut[0186] =  9'sd226;
	icos_lut[0186] = -9'sd94;
	qsin_lut[0187] =  9'sd204;
	icos_lut[0187] = -9'sd136;
	qsin_lut[0188] =  9'sd173;
	icos_lut[0188] = -9'sd173;
	qsin_lut[0189] =  9'sd136;
	icos_lut[0189] = -9'sd204;
	qsin_lut[0190] =  9'sd94;
	icos_lut[0190] = -9'sd226;
	qsin_lut[0191] =  9'sd48;
	icos_lut[0191] = -9'sd240;
	qsin_lut[0192] =  9'sd0;
	icos_lut[0192] = -9'sd243;
	qsin_lut[0193] = -9'sd47;
	icos_lut[0193] = -9'sd238;
	qsin_lut[0194] = -9'sd93;
	icos_lut[0194] = -9'sd225;
	qsin_lut[0195] = -9'sd135;
	icos_lut[0195] = -9'sd202;
	qsin_lut[0196] = -9'sd172;
	icos_lut[0196] = -9'sd172;
	qsin_lut[0197] = -9'sd202;
	icos_lut[0197] = -9'sd135;
	qsin_lut[0198] = -9'sd225;
	icos_lut[0198] = -9'sd93;
	qsin_lut[0199] = -9'sd238;
	icos_lut[0199] = -9'sd47;
	qsin_lut[0200] = -9'sd243;
	icos_lut[0200] = -9'sd0;
	qsin_lut[0201] = -9'sd238;
	icos_lut[0201] =  9'sd47;
	qsin_lut[0202] = -9'sd225;
	icos_lut[0202] =  9'sd93;
	qsin_lut[0203] = -9'sd202;
	icos_lut[0203] =  9'sd135;
	qsin_lut[0204] = -9'sd172;
	icos_lut[0204] =  9'sd172;
	qsin_lut[0205] = -9'sd135;
	icos_lut[0205] =  9'sd202;
	qsin_lut[0206] = -9'sd93;
	icos_lut[0206] =  9'sd225;
	qsin_lut[0207] = -9'sd47;
	icos_lut[0207] =  9'sd238;
	qsin_lut[0208] = -9'sd0;
	icos_lut[0208] =  9'sd243;
	qsin_lut[0209] =  9'sd47;
	icos_lut[0209] =  9'sd238;
	qsin_lut[0210] =  9'sd93;
	icos_lut[0210] =  9'sd225;
	qsin_lut[0211] =  9'sd135;
	icos_lut[0211] =  9'sd202;
	qsin_lut[0212] =  9'sd172;
	icos_lut[0212] =  9'sd172;
	qsin_lut[0213] =  9'sd202;
	icos_lut[0213] =  9'sd135;
	qsin_lut[0214] =  9'sd225;
	icos_lut[0214] =  9'sd93;
	qsin_lut[0215] =  9'sd238;
	icos_lut[0215] =  9'sd47;
	qsin_lut[0216] =  9'sd243;
	icos_lut[0216] =  9'sd0;
	qsin_lut[0217] =  9'sd238;
	icos_lut[0217] = -9'sd47;
	qsin_lut[0218] =  9'sd225;
	icos_lut[0218] = -9'sd93;
	qsin_lut[0219] =  9'sd202;
	icos_lut[0219] = -9'sd135;
	qsin_lut[0220] =  9'sd172;
	icos_lut[0220] = -9'sd172;
	qsin_lut[0221] =  9'sd135;
	icos_lut[0221] = -9'sd202;
	qsin_lut[0222] =  9'sd93;
	icos_lut[0222] = -9'sd225;
	qsin_lut[0223] =  9'sd47;
	icos_lut[0223] = -9'sd238;
	qsin_lut[0224] =  9'sd0;
	icos_lut[0224] = -9'sd241;
	qsin_lut[0225] = -9'sd47;
	icos_lut[0225] = -9'sd236;
	qsin_lut[0226] = -9'sd92;
	icos_lut[0226] = -9'sd223;
	qsin_lut[0227] = -9'sd134;
	icos_lut[0227] = -9'sd200;
	qsin_lut[0228] = -9'sd170;
	icos_lut[0228] = -9'sd170;
	qsin_lut[0229] = -9'sd200;
	icos_lut[0229] = -9'sd134;
	qsin_lut[0230] = -9'sd223;
	icos_lut[0230] = -9'sd92;
	qsin_lut[0231] = -9'sd236;
	icos_lut[0231] = -9'sd47;
	qsin_lut[0232] = -9'sd241;
	icos_lut[0232] = -9'sd0;
	qsin_lut[0233] = -9'sd236;
	icos_lut[0233] =  9'sd47;
	qsin_lut[0234] = -9'sd223;
	icos_lut[0234] =  9'sd92;
	qsin_lut[0235] = -9'sd200;
	icos_lut[0235] =  9'sd134;
	qsin_lut[0236] = -9'sd170;
	icos_lut[0236] =  9'sd170;
	qsin_lut[0237] = -9'sd134;
	icos_lut[0237] =  9'sd200;
	qsin_lut[0238] = -9'sd92;
	icos_lut[0238] =  9'sd223;
	qsin_lut[0239] = -9'sd47;
	icos_lut[0239] =  9'sd236;
	qsin_lut[0240] = -9'sd0;
	icos_lut[0240] =  9'sd241;
	qsin_lut[0241] =  9'sd47;
	icos_lut[0241] =  9'sd236;
	qsin_lut[0242] =  9'sd92;
	icos_lut[0242] =  9'sd223;
	qsin_lut[0243] =  9'sd134;
	icos_lut[0243] =  9'sd200;
	qsin_lut[0244] =  9'sd170;
	icos_lut[0244] =  9'sd170;
	qsin_lut[0245] =  9'sd200;
	icos_lut[0245] =  9'sd134;
	qsin_lut[0246] =  9'sd223;
	icos_lut[0246] =  9'sd92;
	qsin_lut[0247] =  9'sd236;
	icos_lut[0247] =  9'sd47;
	qsin_lut[0248] =  9'sd241;
	icos_lut[0248] =  9'sd0;
	qsin_lut[0249] =  9'sd236;
	icos_lut[0249] = -9'sd47;
	qsin_lut[0250] =  9'sd223;
	icos_lut[0250] = -9'sd92;
	qsin_lut[0251] =  9'sd200;
	icos_lut[0251] = -9'sd134;
	qsin_lut[0252] =  9'sd170;
	icos_lut[0252] = -9'sd170;
	qsin_lut[0253] =  9'sd134;
	icos_lut[0253] = -9'sd200;
	qsin_lut[0254] =  9'sd92;
	icos_lut[0254] = -9'sd223;
	qsin_lut[0255] =  9'sd47;
	icos_lut[0255] = -9'sd236;
	qsin_lut[0256] =  9'sd0;
	icos_lut[0256] = -9'sd239;
	qsin_lut[0257] = -9'sd47;
	icos_lut[0257] = -9'sd234;
	qsin_lut[0258] = -9'sd91;
	icos_lut[0258] = -9'sd221;
	qsin_lut[0259] = -9'sd133;
	icos_lut[0259] = -9'sd199;
	qsin_lut[0260] = -9'sd169;
	icos_lut[0260] = -9'sd169;
	qsin_lut[0261] = -9'sd199;
	icos_lut[0261] = -9'sd133;
	qsin_lut[0262] = -9'sd221;
	icos_lut[0262] = -9'sd91;
	qsin_lut[0263] = -9'sd234;
	icos_lut[0263] = -9'sd47;
	qsin_lut[0264] = -9'sd239;
	icos_lut[0264] = -9'sd0;
	qsin_lut[0265] = -9'sd234;
	icos_lut[0265] =  9'sd47;
	qsin_lut[0266] = -9'sd221;
	icos_lut[0266] =  9'sd91;
	qsin_lut[0267] = -9'sd199;
	icos_lut[0267] =  9'sd133;
	qsin_lut[0268] = -9'sd169;
	icos_lut[0268] =  9'sd169;
	qsin_lut[0269] = -9'sd133;
	icos_lut[0269] =  9'sd199;
	qsin_lut[0270] = -9'sd91;
	icos_lut[0270] =  9'sd221;
	qsin_lut[0271] = -9'sd47;
	icos_lut[0271] =  9'sd234;
	qsin_lut[0272] = -9'sd0;
	icos_lut[0272] =  9'sd239;
	qsin_lut[0273] =  9'sd47;
	icos_lut[0273] =  9'sd234;
	qsin_lut[0274] =  9'sd91;
	icos_lut[0274] =  9'sd221;
	qsin_lut[0275] =  9'sd133;
	icos_lut[0275] =  9'sd199;
	qsin_lut[0276] =  9'sd169;
	icos_lut[0276] =  9'sd169;
	qsin_lut[0277] =  9'sd199;
	icos_lut[0277] =  9'sd133;
	qsin_lut[0278] =  9'sd221;
	icos_lut[0278] =  9'sd91;
	qsin_lut[0279] =  9'sd234;
	icos_lut[0279] =  9'sd47;
	qsin_lut[0280] =  9'sd239;
	icos_lut[0280] =  9'sd0;
	qsin_lut[0281] =  9'sd234;
	icos_lut[0281] = -9'sd47;
	qsin_lut[0282] =  9'sd221;
	icos_lut[0282] = -9'sd91;
	qsin_lut[0283] =  9'sd199;
	icos_lut[0283] = -9'sd133;
	qsin_lut[0284] =  9'sd169;
	icos_lut[0284] = -9'sd169;
	qsin_lut[0285] =  9'sd133;
	icos_lut[0285] = -9'sd199;
	qsin_lut[0286] =  9'sd91;
	icos_lut[0286] = -9'sd221;
	qsin_lut[0287] =  9'sd47;
	icos_lut[0287] = -9'sd234;
	qsin_lut[0288] =  9'sd0;
	icos_lut[0288] = -9'sd237;
	qsin_lut[0289] = -9'sd46;
	icos_lut[0289] = -9'sd232;
	qsin_lut[0290] = -9'sd91;
	icos_lut[0290] = -9'sd219;
	qsin_lut[0291] = -9'sd132;
	icos_lut[0291] = -9'sd197;
	qsin_lut[0292] = -9'sd168;
	icos_lut[0292] = -9'sd168;
	qsin_lut[0293] = -9'sd197;
	icos_lut[0293] = -9'sd132;
	qsin_lut[0294] = -9'sd219;
	icos_lut[0294] = -9'sd91;
	qsin_lut[0295] = -9'sd232;
	icos_lut[0295] = -9'sd46;
	qsin_lut[0296] = -9'sd237;
	icos_lut[0296] = -9'sd0;
	qsin_lut[0297] = -9'sd232;
	icos_lut[0297] =  9'sd46;
	qsin_lut[0298] = -9'sd219;
	icos_lut[0298] =  9'sd91;
	qsin_lut[0299] = -9'sd197;
	icos_lut[0299] =  9'sd132;
	qsin_lut[0300] = -9'sd168;
	icos_lut[0300] =  9'sd168;
	qsin_lut[0301] = -9'sd132;
	icos_lut[0301] =  9'sd197;
	qsin_lut[0302] = -9'sd91;
	icos_lut[0302] =  9'sd219;
	qsin_lut[0303] = -9'sd46;
	icos_lut[0303] =  9'sd232;
	qsin_lut[0304] = -9'sd0;
	icos_lut[0304] =  9'sd237;
	qsin_lut[0305] =  9'sd46;
	icos_lut[0305] =  9'sd232;
	qsin_lut[0306] =  9'sd91;
	icos_lut[0306] =  9'sd219;
	qsin_lut[0307] =  9'sd132;
	icos_lut[0307] =  9'sd197;
	qsin_lut[0308] =  9'sd168;
	icos_lut[0308] =  9'sd168;
	qsin_lut[0309] =  9'sd197;
	icos_lut[0309] =  9'sd132;
	qsin_lut[0310] =  9'sd219;
	icos_lut[0310] =  9'sd91;
	qsin_lut[0311] =  9'sd232;
	icos_lut[0311] =  9'sd46;
	qsin_lut[0312] =  9'sd237;
	icos_lut[0312] =  9'sd0;
	qsin_lut[0313] =  9'sd232;
	icos_lut[0313] = -9'sd46;
	qsin_lut[0314] =  9'sd219;
	icos_lut[0314] = -9'sd91;
	qsin_lut[0315] =  9'sd197;
	icos_lut[0315] = -9'sd132;
	qsin_lut[0316] =  9'sd168;
	icos_lut[0316] = -9'sd168;
	qsin_lut[0317] =  9'sd132;
	icos_lut[0317] = -9'sd197;
	qsin_lut[0318] =  9'sd91;
	icos_lut[0318] = -9'sd219;
	qsin_lut[0319] =  9'sd46;
	icos_lut[0319] = -9'sd232;
	qsin_lut[0320] =  9'sd0;
	icos_lut[0320] = -9'sd235;
	qsin_lut[0321] = -9'sd46;
	icos_lut[0321] = -9'sd230;
	qsin_lut[0322] = -9'sd90;
	icos_lut[0322] = -9'sd217;
	qsin_lut[0323] = -9'sd131;
	icos_lut[0323] = -9'sd195;
	qsin_lut[0324] = -9'sd166;
	icos_lut[0324] = -9'sd166;
	qsin_lut[0325] = -9'sd195;
	icos_lut[0325] = -9'sd131;
	qsin_lut[0326] = -9'sd217;
	icos_lut[0326] = -9'sd90;
	qsin_lut[0327] = -9'sd230;
	icos_lut[0327] = -9'sd46;
	qsin_lut[0328] = -9'sd235;
	icos_lut[0328] = -9'sd0;
	qsin_lut[0329] = -9'sd230;
	icos_lut[0329] =  9'sd46;
	qsin_lut[0330] = -9'sd217;
	icos_lut[0330] =  9'sd90;
	qsin_lut[0331] = -9'sd195;
	icos_lut[0331] =  9'sd131;
	qsin_lut[0332] = -9'sd166;
	icos_lut[0332] =  9'sd166;
	qsin_lut[0333] = -9'sd131;
	icos_lut[0333] =  9'sd195;
	qsin_lut[0334] = -9'sd90;
	icos_lut[0334] =  9'sd217;
	qsin_lut[0335] = -9'sd46;
	icos_lut[0335] =  9'sd230;
	qsin_lut[0336] = -9'sd0;
	icos_lut[0336] =  9'sd235;
	qsin_lut[0337] =  9'sd46;
	icos_lut[0337] =  9'sd230;
	qsin_lut[0338] =  9'sd90;
	icos_lut[0338] =  9'sd217;
	qsin_lut[0339] =  9'sd131;
	icos_lut[0339] =  9'sd195;
	qsin_lut[0340] =  9'sd166;
	icos_lut[0340] =  9'sd166;
	qsin_lut[0341] =  9'sd195;
	icos_lut[0341] =  9'sd131;
	qsin_lut[0342] =  9'sd217;
	icos_lut[0342] =  9'sd90;
	qsin_lut[0343] =  9'sd230;
	icos_lut[0343] =  9'sd46;
	qsin_lut[0344] =  9'sd235;
	icos_lut[0344] =  9'sd0;
	qsin_lut[0345] =  9'sd230;
	icos_lut[0345] = -9'sd46;
	qsin_lut[0346] =  9'sd217;
	icos_lut[0346] = -9'sd90;
	qsin_lut[0347] =  9'sd195;
	icos_lut[0347] = -9'sd131;
	qsin_lut[0348] =  9'sd166;
	icos_lut[0348] = -9'sd166;
	qsin_lut[0349] =  9'sd131;
	icos_lut[0349] = -9'sd195;
	qsin_lut[0350] =  9'sd90;
	icos_lut[0350] = -9'sd217;
	qsin_lut[0351] =  9'sd46;
	icos_lut[0351] = -9'sd230;
	qsin_lut[0352] =  9'sd0;
	icos_lut[0352] = -9'sd233;
	qsin_lut[0353] = -9'sd45;
	icos_lut[0353] = -9'sd229;
	qsin_lut[0354] = -9'sd89;
	icos_lut[0354] = -9'sd215;
	qsin_lut[0355] = -9'sd129;
	icos_lut[0355] = -9'sd194;
	qsin_lut[0356] = -9'sd165;
	icos_lut[0356] = -9'sd165;
	qsin_lut[0357] = -9'sd194;
	icos_lut[0357] = -9'sd129;
	qsin_lut[0358] = -9'sd215;
	icos_lut[0358] = -9'sd89;
	qsin_lut[0359] = -9'sd229;
	icos_lut[0359] = -9'sd45;
	qsin_lut[0360] = -9'sd233;
	icos_lut[0360] = -9'sd0;
	qsin_lut[0361] = -9'sd229;
	icos_lut[0361] =  9'sd45;
	qsin_lut[0362] = -9'sd215;
	icos_lut[0362] =  9'sd89;
	qsin_lut[0363] = -9'sd194;
	icos_lut[0363] =  9'sd129;
	qsin_lut[0364] = -9'sd165;
	icos_lut[0364] =  9'sd165;
	qsin_lut[0365] = -9'sd129;
	icos_lut[0365] =  9'sd194;
	qsin_lut[0366] = -9'sd89;
	icos_lut[0366] =  9'sd215;
	qsin_lut[0367] = -9'sd45;
	icos_lut[0367] =  9'sd229;
	qsin_lut[0368] = -9'sd0;
	icos_lut[0368] =  9'sd233;
	qsin_lut[0369] =  9'sd45;
	icos_lut[0369] =  9'sd229;
	qsin_lut[0370] =  9'sd89;
	icos_lut[0370] =  9'sd215;
	qsin_lut[0371] =  9'sd129;
	icos_lut[0371] =  9'sd194;
	qsin_lut[0372] =  9'sd165;
	icos_lut[0372] =  9'sd165;
	qsin_lut[0373] =  9'sd194;
	icos_lut[0373] =  9'sd129;
	qsin_lut[0374] =  9'sd215;
	icos_lut[0374] =  9'sd89;
	qsin_lut[0375] =  9'sd229;
	icos_lut[0375] =  9'sd45;
	qsin_lut[0376] =  9'sd233;
	icos_lut[0376] =  9'sd0;
	qsin_lut[0377] =  9'sd229;
	icos_lut[0377] = -9'sd45;
	qsin_lut[0378] =  9'sd215;
	icos_lut[0378] = -9'sd89;
	qsin_lut[0379] =  9'sd194;
	icos_lut[0379] = -9'sd129;
	qsin_lut[0380] =  9'sd165;
	icos_lut[0380] = -9'sd165;
	qsin_lut[0381] =  9'sd129;
	icos_lut[0381] = -9'sd194;
	qsin_lut[0382] =  9'sd89;
	icos_lut[0382] = -9'sd215;
	qsin_lut[0383] =  9'sd45;
	icos_lut[0383] = -9'sd229;
	qsin_lut[0384] =  9'sd0;
	icos_lut[0384] = -9'sd231;
	qsin_lut[0385] = -9'sd45;
	icos_lut[0385] = -9'sd227;
	qsin_lut[0386] = -9'sd88;
	icos_lut[0386] = -9'sd213;
	qsin_lut[0387] = -9'sd128;
	icos_lut[0387] = -9'sd192;
	qsin_lut[0388] = -9'sd163;
	icos_lut[0388] = -9'sd163;
	qsin_lut[0389] = -9'sd192;
	icos_lut[0389] = -9'sd128;
	qsin_lut[0390] = -9'sd213;
	icos_lut[0390] = -9'sd88;
	qsin_lut[0391] = -9'sd227;
	icos_lut[0391] = -9'sd45;
	qsin_lut[0392] = -9'sd231;
	icos_lut[0392] = -9'sd0;
	qsin_lut[0393] = -9'sd227;
	icos_lut[0393] =  9'sd45;
	qsin_lut[0394] = -9'sd213;
	icos_lut[0394] =  9'sd88;
	qsin_lut[0395] = -9'sd192;
	icos_lut[0395] =  9'sd128;
	qsin_lut[0396] = -9'sd163;
	icos_lut[0396] =  9'sd163;
	qsin_lut[0397] = -9'sd128;
	icos_lut[0397] =  9'sd192;
	qsin_lut[0398] = -9'sd88;
	icos_lut[0398] =  9'sd213;
	qsin_lut[0399] = -9'sd45;
	icos_lut[0399] =  9'sd227;
	qsin_lut[0400] = -9'sd0;
	icos_lut[0400] =  9'sd231;
	qsin_lut[0401] =  9'sd45;
	icos_lut[0401] =  9'sd227;
	qsin_lut[0402] =  9'sd88;
	icos_lut[0402] =  9'sd213;
	qsin_lut[0403] =  9'sd128;
	icos_lut[0403] =  9'sd192;
	qsin_lut[0404] =  9'sd163;
	icos_lut[0404] =  9'sd163;
	qsin_lut[0405] =  9'sd192;
	icos_lut[0405] =  9'sd128;
	qsin_lut[0406] =  9'sd213;
	icos_lut[0406] =  9'sd88;
	qsin_lut[0407] =  9'sd227;
	icos_lut[0407] =  9'sd45;
	qsin_lut[0408] =  9'sd231;
	icos_lut[0408] =  9'sd0;
	qsin_lut[0409] =  9'sd227;
	icos_lut[0409] = -9'sd45;
	qsin_lut[0410] =  9'sd213;
	icos_lut[0410] = -9'sd88;
	qsin_lut[0411] =  9'sd192;
	icos_lut[0411] = -9'sd128;
	qsin_lut[0412] =  9'sd163;
	icos_lut[0412] = -9'sd163;
	qsin_lut[0413] =  9'sd128;
	icos_lut[0413] = -9'sd192;
	qsin_lut[0414] =  9'sd88;
	icos_lut[0414] = -9'sd213;
	qsin_lut[0415] =  9'sd45;
	icos_lut[0415] = -9'sd227;
	qsin_lut[0416] =  9'sd0;
	icos_lut[0416] = -9'sd229;
	qsin_lut[0417] = -9'sd45;
	icos_lut[0417] = -9'sd225;
	qsin_lut[0418] = -9'sd88;
	icos_lut[0418] = -9'sd212;
	qsin_lut[0419] = -9'sd127;
	icos_lut[0419] = -9'sd190;
	qsin_lut[0420] = -9'sd162;
	icos_lut[0420] = -9'sd162;
	qsin_lut[0421] = -9'sd190;
	icos_lut[0421] = -9'sd127;
	qsin_lut[0422] = -9'sd212;
	icos_lut[0422] = -9'sd88;
	qsin_lut[0423] = -9'sd225;
	icos_lut[0423] = -9'sd45;
	qsin_lut[0424] = -9'sd229;
	icos_lut[0424] = -9'sd0;
	qsin_lut[0425] = -9'sd225;
	icos_lut[0425] =  9'sd45;
	qsin_lut[0426] = -9'sd212;
	icos_lut[0426] =  9'sd88;
	qsin_lut[0427] = -9'sd190;
	icos_lut[0427] =  9'sd127;
	qsin_lut[0428] = -9'sd162;
	icos_lut[0428] =  9'sd162;
	qsin_lut[0429] = -9'sd127;
	icos_lut[0429] =  9'sd190;
	qsin_lut[0430] = -9'sd88;
	icos_lut[0430] =  9'sd212;
	qsin_lut[0431] = -9'sd45;
	icos_lut[0431] =  9'sd225;
	qsin_lut[0432] = -9'sd0;
	icos_lut[0432] =  9'sd229;
	qsin_lut[0433] =  9'sd45;
	icos_lut[0433] =  9'sd225;
	qsin_lut[0434] =  9'sd88;
	icos_lut[0434] =  9'sd212;
	qsin_lut[0435] =  9'sd127;
	icos_lut[0435] =  9'sd190;
	qsin_lut[0436] =  9'sd162;
	icos_lut[0436] =  9'sd162;
	qsin_lut[0437] =  9'sd190;
	icos_lut[0437] =  9'sd127;
	qsin_lut[0438] =  9'sd212;
	icos_lut[0438] =  9'sd88;
	qsin_lut[0439] =  9'sd225;
	icos_lut[0439] =  9'sd45;
	qsin_lut[0440] =  9'sd229;
	icos_lut[0440] =  9'sd0;
	qsin_lut[0441] =  9'sd225;
	icos_lut[0441] = -9'sd45;
	qsin_lut[0442] =  9'sd212;
	icos_lut[0442] = -9'sd88;
	qsin_lut[0443] =  9'sd190;
	icos_lut[0443] = -9'sd127;
	qsin_lut[0444] =  9'sd162;
	icos_lut[0444] = -9'sd162;
	qsin_lut[0445] =  9'sd127;
	icos_lut[0445] = -9'sd190;
	qsin_lut[0446] =  9'sd88;
	icos_lut[0446] = -9'sd212;
	qsin_lut[0447] =  9'sd45;
	icos_lut[0447] = -9'sd225;
	qsin_lut[0448] =  9'sd0;
	icos_lut[0448] = -9'sd227;
	qsin_lut[0449] = -9'sd44;
	icos_lut[0449] = -9'sd223;
	qsin_lut[0450] = -9'sd87;
	icos_lut[0450] = -9'sd210;
	qsin_lut[0451] = -9'sd126;
	icos_lut[0451] = -9'sd189;
	qsin_lut[0452] = -9'sd161;
	icos_lut[0452] = -9'sd161;
	qsin_lut[0453] = -9'sd189;
	icos_lut[0453] = -9'sd126;
	qsin_lut[0454] = -9'sd210;
	icos_lut[0454] = -9'sd87;
	qsin_lut[0455] = -9'sd223;
	icos_lut[0455] = -9'sd44;
	qsin_lut[0456] = -9'sd227;
	icos_lut[0456] = -9'sd0;
	qsin_lut[0457] = -9'sd223;
	icos_lut[0457] =  9'sd44;
	qsin_lut[0458] = -9'sd210;
	icos_lut[0458] =  9'sd87;
	qsin_lut[0459] = -9'sd189;
	icos_lut[0459] =  9'sd126;
	qsin_lut[0460] = -9'sd161;
	icos_lut[0460] =  9'sd161;
	qsin_lut[0461] = -9'sd126;
	icos_lut[0461] =  9'sd189;
	qsin_lut[0462] = -9'sd87;
	icos_lut[0462] =  9'sd210;
	qsin_lut[0463] = -9'sd44;
	icos_lut[0463] =  9'sd223;
	qsin_lut[0464] = -9'sd0;
	icos_lut[0464] =  9'sd227;
	qsin_lut[0465] =  9'sd44;
	icos_lut[0465] =  9'sd223;
	qsin_lut[0466] =  9'sd87;
	icos_lut[0466] =  9'sd210;
	qsin_lut[0467] =  9'sd126;
	icos_lut[0467] =  9'sd189;
	qsin_lut[0468] =  9'sd161;
	icos_lut[0468] =  9'sd161;
	qsin_lut[0469] =  9'sd189;
	icos_lut[0469] =  9'sd126;
	qsin_lut[0470] =  9'sd210;
	icos_lut[0470] =  9'sd87;
	qsin_lut[0471] =  9'sd223;
	icos_lut[0471] =  9'sd44;
	qsin_lut[0472] =  9'sd227;
	icos_lut[0472] =  9'sd0;
	qsin_lut[0473] =  9'sd223;
	icos_lut[0473] = -9'sd44;
	qsin_lut[0474] =  9'sd210;
	icos_lut[0474] = -9'sd87;
	qsin_lut[0475] =  9'sd189;
	icos_lut[0475] = -9'sd126;
	qsin_lut[0476] =  9'sd161;
	icos_lut[0476] = -9'sd161;
	qsin_lut[0477] =  9'sd126;
	icos_lut[0477] = -9'sd189;
	qsin_lut[0478] =  9'sd87;
	icos_lut[0478] = -9'sd210;
	qsin_lut[0479] =  9'sd44;
	icos_lut[0479] = -9'sd223;
	qsin_lut[0480] =  9'sd0;
	icos_lut[0480] = -9'sd225;
	qsin_lut[0481] = -9'sd44;
	icos_lut[0481] = -9'sd221;
	qsin_lut[0482] = -9'sd86;
	icos_lut[0482] = -9'sd208;
	qsin_lut[0483] = -9'sd125;
	icos_lut[0483] = -9'sd187;
	qsin_lut[0484] = -9'sd159;
	icos_lut[0484] = -9'sd159;
	qsin_lut[0485] = -9'sd187;
	icos_lut[0485] = -9'sd125;
	qsin_lut[0486] = -9'sd208;
	icos_lut[0486] = -9'sd86;
	qsin_lut[0487] = -9'sd221;
	icos_lut[0487] = -9'sd44;
	qsin_lut[0488] = -9'sd225;
	icos_lut[0488] = -9'sd0;
	qsin_lut[0489] = -9'sd221;
	icos_lut[0489] =  9'sd44;
	qsin_lut[0490] = -9'sd208;
	icos_lut[0490] =  9'sd86;
	qsin_lut[0491] = -9'sd187;
	icos_lut[0491] =  9'sd125;
	qsin_lut[0492] = -9'sd159;
	icos_lut[0492] =  9'sd159;
	qsin_lut[0493] = -9'sd125;
	icos_lut[0493] =  9'sd187;
	qsin_lut[0494] = -9'sd86;
	icos_lut[0494] =  9'sd208;
	qsin_lut[0495] = -9'sd44;
	icos_lut[0495] =  9'sd221;
	qsin_lut[0496] = -9'sd0;
	icos_lut[0496] =  9'sd225;
	qsin_lut[0497] =  9'sd44;
	icos_lut[0497] =  9'sd221;
	qsin_lut[0498] =  9'sd86;
	icos_lut[0498] =  9'sd208;
	qsin_lut[0499] =  9'sd125;
	icos_lut[0499] =  9'sd187;
	qsin_lut[0500] =  9'sd159;
	icos_lut[0500] =  9'sd159;
	qsin_lut[0501] =  9'sd187;
	icos_lut[0501] =  9'sd125;
	qsin_lut[0502] =  9'sd208;
	icos_lut[0502] =  9'sd86;
	qsin_lut[0503] =  9'sd221;
	icos_lut[0503] =  9'sd44;
	qsin_lut[0504] =  9'sd225;
	icos_lut[0504] =  9'sd0;
	qsin_lut[0505] =  9'sd221;
	icos_lut[0505] = -9'sd44;
	qsin_lut[0506] =  9'sd208;
	icos_lut[0506] = -9'sd86;
	qsin_lut[0507] =  9'sd187;
	icos_lut[0507] = -9'sd125;
	qsin_lut[0508] =  9'sd159;
	icos_lut[0508] = -9'sd159;
	qsin_lut[0509] =  9'sd125;
	icos_lut[0509] = -9'sd187;
	qsin_lut[0510] =  9'sd86;
	icos_lut[0510] = -9'sd208;
	qsin_lut[0511] =  9'sd44;
	icos_lut[0511] = -9'sd221;
	qsin_lut[0512] =  9'sd0;
	icos_lut[0512] = -9'sd223;
	qsin_lut[0513] = -9'sd44;
	icos_lut[0513] = -9'sd219;
	qsin_lut[0514] = -9'sd85;
	icos_lut[0514] = -9'sd206;
	qsin_lut[0515] = -9'sd124;
	icos_lut[0515] = -9'sd185;
	qsin_lut[0516] = -9'sd158;
	icos_lut[0516] = -9'sd158;
	qsin_lut[0517] = -9'sd185;
	icos_lut[0517] = -9'sd124;
	qsin_lut[0518] = -9'sd206;
	icos_lut[0518] = -9'sd85;
	qsin_lut[0519] = -9'sd219;
	icos_lut[0519] = -9'sd44;
	qsin_lut[0520] = -9'sd223;
	icos_lut[0520] = -9'sd0;
	qsin_lut[0521] = -9'sd219;
	icos_lut[0521] =  9'sd44;
	qsin_lut[0522] = -9'sd206;
	icos_lut[0522] =  9'sd85;
	qsin_lut[0523] = -9'sd185;
	icos_lut[0523] =  9'sd124;
	qsin_lut[0524] = -9'sd158;
	icos_lut[0524] =  9'sd158;
	qsin_lut[0525] = -9'sd124;
	icos_lut[0525] =  9'sd185;
	qsin_lut[0526] = -9'sd85;
	icos_lut[0526] =  9'sd206;
	qsin_lut[0527] = -9'sd44;
	icos_lut[0527] =  9'sd219;
	qsin_lut[0528] = -9'sd0;
	icos_lut[0528] =  9'sd223;
	qsin_lut[0529] =  9'sd44;
	icos_lut[0529] =  9'sd219;
	qsin_lut[0530] =  9'sd85;
	icos_lut[0530] =  9'sd206;
	qsin_lut[0531] =  9'sd124;
	icos_lut[0531] =  9'sd185;
	qsin_lut[0532] =  9'sd158;
	icos_lut[0532] =  9'sd158;
	qsin_lut[0533] =  9'sd185;
	icos_lut[0533] =  9'sd124;
	qsin_lut[0534] =  9'sd206;
	icos_lut[0534] =  9'sd85;
	qsin_lut[0535] =  9'sd219;
	icos_lut[0535] =  9'sd44;
	qsin_lut[0536] =  9'sd223;
	icos_lut[0536] =  9'sd0;
	qsin_lut[0537] =  9'sd219;
	icos_lut[0537] = -9'sd44;
	qsin_lut[0538] =  9'sd206;
	icos_lut[0538] = -9'sd85;
	qsin_lut[0539] =  9'sd185;
	icos_lut[0539] = -9'sd124;
	qsin_lut[0540] =  9'sd158;
	icos_lut[0540] = -9'sd158;
	qsin_lut[0541] =  9'sd124;
	icos_lut[0541] = -9'sd185;
	qsin_lut[0542] =  9'sd85;
	icos_lut[0542] = -9'sd206;
	qsin_lut[0543] =  9'sd44;
	icos_lut[0543] = -9'sd219;
	qsin_lut[0544] =  9'sd0;
	icos_lut[0544] = -9'sd221;
	qsin_lut[0545] = -9'sd43;
	icos_lut[0545] = -9'sd217;
	qsin_lut[0546] = -9'sd85;
	icos_lut[0546] = -9'sd204;
	qsin_lut[0547] = -9'sd123;
	icos_lut[0547] = -9'sd184;
	qsin_lut[0548] = -9'sd156;
	icos_lut[0548] = -9'sd156;
	qsin_lut[0549] = -9'sd184;
	icos_lut[0549] = -9'sd123;
	qsin_lut[0550] = -9'sd204;
	icos_lut[0550] = -9'sd85;
	qsin_lut[0551] = -9'sd217;
	icos_lut[0551] = -9'sd43;
	qsin_lut[0552] = -9'sd221;
	icos_lut[0552] = -9'sd0;
	qsin_lut[0553] = -9'sd217;
	icos_lut[0553] =  9'sd43;
	qsin_lut[0554] = -9'sd204;
	icos_lut[0554] =  9'sd85;
	qsin_lut[0555] = -9'sd184;
	icos_lut[0555] =  9'sd123;
	qsin_lut[0556] = -9'sd156;
	icos_lut[0556] =  9'sd156;
	qsin_lut[0557] = -9'sd123;
	icos_lut[0557] =  9'sd184;
	qsin_lut[0558] = -9'sd85;
	icos_lut[0558] =  9'sd204;
	qsin_lut[0559] = -9'sd43;
	icos_lut[0559] =  9'sd217;
	qsin_lut[0560] = -9'sd0;
	icos_lut[0560] =  9'sd221;
	qsin_lut[0561] =  9'sd43;
	icos_lut[0561] =  9'sd217;
	qsin_lut[0562] =  9'sd85;
	icos_lut[0562] =  9'sd204;
	qsin_lut[0563] =  9'sd123;
	icos_lut[0563] =  9'sd184;
	qsin_lut[0564] =  9'sd156;
	icos_lut[0564] =  9'sd156;
	qsin_lut[0565] =  9'sd184;
	icos_lut[0565] =  9'sd123;
	qsin_lut[0566] =  9'sd204;
	icos_lut[0566] =  9'sd85;
	qsin_lut[0567] =  9'sd217;
	icos_lut[0567] =  9'sd43;
	qsin_lut[0568] =  9'sd221;
	icos_lut[0568] =  9'sd0;
	qsin_lut[0569] =  9'sd217;
	icos_lut[0569] = -9'sd43;
	qsin_lut[0570] =  9'sd204;
	icos_lut[0570] = -9'sd85;
	qsin_lut[0571] =  9'sd184;
	icos_lut[0571] = -9'sd123;
	qsin_lut[0572] =  9'sd156;
	icos_lut[0572] = -9'sd156;
	qsin_lut[0573] =  9'sd123;
	icos_lut[0573] = -9'sd184;
	qsin_lut[0574] =  9'sd85;
	icos_lut[0574] = -9'sd204;
	qsin_lut[0575] =  9'sd43;
	icos_lut[0575] = -9'sd217;
	qsin_lut[0576] =  9'sd0;
	icos_lut[0576] = -9'sd219;
	qsin_lut[0577] = -9'sd43;
	icos_lut[0577] = -9'sd215;
	qsin_lut[0578] = -9'sd84;
	icos_lut[0578] = -9'sd202;
	qsin_lut[0579] = -9'sd122;
	icos_lut[0579] = -9'sd182;
	qsin_lut[0580] = -9'sd155;
	icos_lut[0580] = -9'sd155;
	qsin_lut[0581] = -9'sd182;
	icos_lut[0581] = -9'sd122;
	qsin_lut[0582] = -9'sd202;
	icos_lut[0582] = -9'sd84;
	qsin_lut[0583] = -9'sd215;
	icos_lut[0583] = -9'sd43;
	qsin_lut[0584] = -9'sd219;
	icos_lut[0584] = -9'sd0;
	qsin_lut[0585] = -9'sd215;
	icos_lut[0585] =  9'sd43;
	qsin_lut[0586] = -9'sd202;
	icos_lut[0586] =  9'sd84;
	qsin_lut[0587] = -9'sd182;
	icos_lut[0587] =  9'sd122;
	qsin_lut[0588] = -9'sd155;
	icos_lut[0588] =  9'sd155;
	qsin_lut[0589] = -9'sd122;
	icos_lut[0589] =  9'sd182;
	qsin_lut[0590] = -9'sd84;
	icos_lut[0590] =  9'sd202;
	qsin_lut[0591] = -9'sd43;
	icos_lut[0591] =  9'sd215;
	qsin_lut[0592] = -9'sd0;
	icos_lut[0592] =  9'sd219;
	qsin_lut[0593] =  9'sd43;
	icos_lut[0593] =  9'sd215;
	qsin_lut[0594] =  9'sd84;
	icos_lut[0594] =  9'sd202;
	qsin_lut[0595] =  9'sd122;
	icos_lut[0595] =  9'sd182;
	qsin_lut[0596] =  9'sd155;
	icos_lut[0596] =  9'sd155;
	qsin_lut[0597] =  9'sd182;
	icos_lut[0597] =  9'sd122;
	qsin_lut[0598] =  9'sd202;
	icos_lut[0598] =  9'sd84;
	qsin_lut[0599] =  9'sd215;
	icos_lut[0599] =  9'sd43;
	qsin_lut[0600] =  9'sd219;
	icos_lut[0600] =  9'sd0;
	qsin_lut[0601] =  9'sd215;
	icos_lut[0601] = -9'sd43;
	qsin_lut[0602] =  9'sd202;
	icos_lut[0602] = -9'sd84;
	qsin_lut[0603] =  9'sd182;
	icos_lut[0603] = -9'sd122;
	qsin_lut[0604] =  9'sd155;
	icos_lut[0604] = -9'sd155;
	qsin_lut[0605] =  9'sd122;
	icos_lut[0605] = -9'sd182;
	qsin_lut[0606] =  9'sd84;
	icos_lut[0606] = -9'sd202;
	qsin_lut[0607] =  9'sd43;
	icos_lut[0607] = -9'sd215;
	qsin_lut[0608] =  9'sd0;
	icos_lut[0608] = -9'sd217;
	qsin_lut[0609] = -9'sd42;
	icos_lut[0609] = -9'sd213;
	qsin_lut[0610] = -9'sd83;
	icos_lut[0610] = -9'sd200;
	qsin_lut[0611] = -9'sd121;
	icos_lut[0611] = -9'sd180;
	qsin_lut[0612] = -9'sd153;
	icos_lut[0612] = -9'sd153;
	qsin_lut[0613] = -9'sd180;
	icos_lut[0613] = -9'sd121;
	qsin_lut[0614] = -9'sd200;
	icos_lut[0614] = -9'sd83;
	qsin_lut[0615] = -9'sd213;
	icos_lut[0615] = -9'sd42;
	qsin_lut[0616] = -9'sd217;
	icos_lut[0616] = -9'sd0;
	qsin_lut[0617] = -9'sd213;
	icos_lut[0617] =  9'sd42;
	qsin_lut[0618] = -9'sd200;
	icos_lut[0618] =  9'sd83;
	qsin_lut[0619] = -9'sd180;
	icos_lut[0619] =  9'sd121;
	qsin_lut[0620] = -9'sd153;
	icos_lut[0620] =  9'sd153;
	qsin_lut[0621] = -9'sd121;
	icos_lut[0621] =  9'sd180;
	qsin_lut[0622] = -9'sd83;
	icos_lut[0622] =  9'sd200;
	qsin_lut[0623] = -9'sd42;
	icos_lut[0623] =  9'sd213;
	qsin_lut[0624] = -9'sd0;
	icos_lut[0624] =  9'sd217;
	qsin_lut[0625] =  9'sd42;
	icos_lut[0625] =  9'sd213;
	qsin_lut[0626] =  9'sd83;
	icos_lut[0626] =  9'sd200;
	qsin_lut[0627] =  9'sd121;
	icos_lut[0627] =  9'sd180;
	qsin_lut[0628] =  9'sd153;
	icos_lut[0628] =  9'sd153;
	qsin_lut[0629] =  9'sd180;
	icos_lut[0629] =  9'sd121;
	qsin_lut[0630] =  9'sd200;
	icos_lut[0630] =  9'sd83;
	qsin_lut[0631] =  9'sd213;
	icos_lut[0631] =  9'sd42;
	qsin_lut[0632] =  9'sd217;
	icos_lut[0632] =  9'sd0;
	qsin_lut[0633] =  9'sd213;
	icos_lut[0633] = -9'sd42;
	qsin_lut[0634] =  9'sd200;
	icos_lut[0634] = -9'sd83;
	qsin_lut[0635] =  9'sd180;
	icos_lut[0635] = -9'sd121;
	qsin_lut[0636] =  9'sd153;
	icos_lut[0636] = -9'sd153;
	qsin_lut[0637] =  9'sd121;
	icos_lut[0637] = -9'sd180;
	qsin_lut[0638] =  9'sd83;
	icos_lut[0638] = -9'sd200;
	qsin_lut[0639] =  9'sd42;
	icos_lut[0639] = -9'sd213;
	qsin_lut[0640] =  9'sd0;
	icos_lut[0640] = -9'sd215;
	qsin_lut[0641] = -9'sd42;
	icos_lut[0641] = -9'sd211;
	qsin_lut[0642] = -9'sd82;
	icos_lut[0642] = -9'sd199;
	qsin_lut[0643] = -9'sd119;
	icos_lut[0643] = -9'sd179;
	qsin_lut[0644] = -9'sd152;
	icos_lut[0644] = -9'sd152;
	qsin_lut[0645] = -9'sd179;
	icos_lut[0645] = -9'sd119;
	qsin_lut[0646] = -9'sd199;
	icos_lut[0646] = -9'sd82;
	qsin_lut[0647] = -9'sd211;
	icos_lut[0647] = -9'sd42;
	qsin_lut[0648] = -9'sd215;
	icos_lut[0648] = -9'sd0;
	qsin_lut[0649] = -9'sd211;
	icos_lut[0649] =  9'sd42;
	qsin_lut[0650] = -9'sd199;
	icos_lut[0650] =  9'sd82;
	qsin_lut[0651] = -9'sd179;
	icos_lut[0651] =  9'sd119;
	qsin_lut[0652] = -9'sd152;
	icos_lut[0652] =  9'sd152;
	qsin_lut[0653] = -9'sd119;
	icos_lut[0653] =  9'sd179;
	qsin_lut[0654] = -9'sd82;
	icos_lut[0654] =  9'sd199;
	qsin_lut[0655] = -9'sd42;
	icos_lut[0655] =  9'sd211;
	qsin_lut[0656] = -9'sd0;
	icos_lut[0656] =  9'sd215;
	qsin_lut[0657] =  9'sd42;
	icos_lut[0657] =  9'sd211;
	qsin_lut[0658] =  9'sd82;
	icos_lut[0658] =  9'sd199;
	qsin_lut[0659] =  9'sd119;
	icos_lut[0659] =  9'sd179;
	qsin_lut[0660] =  9'sd152;
	icos_lut[0660] =  9'sd152;
	qsin_lut[0661] =  9'sd179;
	icos_lut[0661] =  9'sd119;
	qsin_lut[0662] =  9'sd199;
	icos_lut[0662] =  9'sd82;
	qsin_lut[0663] =  9'sd211;
	icos_lut[0663] =  9'sd42;
	qsin_lut[0664] =  9'sd215;
	icos_lut[0664] =  9'sd0;
	qsin_lut[0665] =  9'sd211;
	icos_lut[0665] = -9'sd42;
	qsin_lut[0666] =  9'sd199;
	icos_lut[0666] = -9'sd82;
	qsin_lut[0667] =  9'sd179;
	icos_lut[0667] = -9'sd119;
	qsin_lut[0668] =  9'sd152;
	icos_lut[0668] = -9'sd152;
	qsin_lut[0669] =  9'sd119;
	icos_lut[0669] = -9'sd179;
	qsin_lut[0670] =  9'sd82;
	icos_lut[0670] = -9'sd199;
	qsin_lut[0671] =  9'sd42;
	icos_lut[0671] = -9'sd211;
	qsin_lut[0672] =  9'sd0;
	icos_lut[0672] = -9'sd213;
	qsin_lut[0673] = -9'sd42;
	icos_lut[0673] = -9'sd209;
	qsin_lut[0674] = -9'sd82;
	icos_lut[0674] = -9'sd197;
	qsin_lut[0675] = -9'sd118;
	icos_lut[0675] = -9'sd177;
	qsin_lut[0676] = -9'sd151;
	icos_lut[0676] = -9'sd151;
	qsin_lut[0677] = -9'sd177;
	icos_lut[0677] = -9'sd118;
	qsin_lut[0678] = -9'sd197;
	icos_lut[0678] = -9'sd82;
	qsin_lut[0679] = -9'sd209;
	icos_lut[0679] = -9'sd42;
	qsin_lut[0680] = -9'sd213;
	icos_lut[0680] = -9'sd0;
	qsin_lut[0681] = -9'sd209;
	icos_lut[0681] =  9'sd42;
	qsin_lut[0682] = -9'sd197;
	icos_lut[0682] =  9'sd82;
	qsin_lut[0683] = -9'sd177;
	icos_lut[0683] =  9'sd118;
	qsin_lut[0684] = -9'sd151;
	icos_lut[0684] =  9'sd151;
	qsin_lut[0685] = -9'sd118;
	icos_lut[0685] =  9'sd177;
	qsin_lut[0686] = -9'sd82;
	icos_lut[0686] =  9'sd197;
	qsin_lut[0687] = -9'sd42;
	icos_lut[0687] =  9'sd209;
	qsin_lut[0688] = -9'sd0;
	icos_lut[0688] =  9'sd213;
	qsin_lut[0689] =  9'sd42;
	icos_lut[0689] =  9'sd209;
	qsin_lut[0690] =  9'sd82;
	icos_lut[0690] =  9'sd197;
	qsin_lut[0691] =  9'sd118;
	icos_lut[0691] =  9'sd177;
	qsin_lut[0692] =  9'sd151;
	icos_lut[0692] =  9'sd151;
	qsin_lut[0693] =  9'sd177;
	icos_lut[0693] =  9'sd118;
	qsin_lut[0694] =  9'sd197;
	icos_lut[0694] =  9'sd82;
	qsin_lut[0695] =  9'sd209;
	icos_lut[0695] =  9'sd42;
	qsin_lut[0696] =  9'sd213;
	icos_lut[0696] =  9'sd0;
	qsin_lut[0697] =  9'sd209;
	icos_lut[0697] = -9'sd42;
	qsin_lut[0698] =  9'sd197;
	icos_lut[0698] = -9'sd82;
	qsin_lut[0699] =  9'sd177;
	icos_lut[0699] = -9'sd118;
	qsin_lut[0700] =  9'sd151;
	icos_lut[0700] = -9'sd151;
	qsin_lut[0701] =  9'sd118;
	icos_lut[0701] = -9'sd177;
	qsin_lut[0702] =  9'sd82;
	icos_lut[0702] = -9'sd197;
	qsin_lut[0703] =  9'sd42;
	icos_lut[0703] = -9'sd209;
	qsin_lut[0704] =  9'sd0;
	icos_lut[0704] = -9'sd211;
	qsin_lut[0705] = -9'sd41;
	icos_lut[0705] = -9'sd207;
	qsin_lut[0706] = -9'sd81;
	icos_lut[0706] = -9'sd195;
	qsin_lut[0707] = -9'sd117;
	icos_lut[0707] = -9'sd175;
	qsin_lut[0708] = -9'sd149;
	icos_lut[0708] = -9'sd149;
	qsin_lut[0709] = -9'sd175;
	icos_lut[0709] = -9'sd117;
	qsin_lut[0710] = -9'sd195;
	icos_lut[0710] = -9'sd81;
	qsin_lut[0711] = -9'sd207;
	icos_lut[0711] = -9'sd41;
	qsin_lut[0712] = -9'sd211;
	icos_lut[0712] = -9'sd0;
	qsin_lut[0713] = -9'sd207;
	icos_lut[0713] =  9'sd41;
	qsin_lut[0714] = -9'sd195;
	icos_lut[0714] =  9'sd81;
	qsin_lut[0715] = -9'sd175;
	icos_lut[0715] =  9'sd117;
	qsin_lut[0716] = -9'sd149;
	icos_lut[0716] =  9'sd149;
	qsin_lut[0717] = -9'sd117;
	icos_lut[0717] =  9'sd175;
	qsin_lut[0718] = -9'sd81;
	icos_lut[0718] =  9'sd195;
	qsin_lut[0719] = -9'sd41;
	icos_lut[0719] =  9'sd207;
	qsin_lut[0720] = -9'sd0;
	icos_lut[0720] =  9'sd211;
	qsin_lut[0721] =  9'sd41;
	icos_lut[0721] =  9'sd207;
	qsin_lut[0722] =  9'sd81;
	icos_lut[0722] =  9'sd195;
	qsin_lut[0723] =  9'sd117;
	icos_lut[0723] =  9'sd175;
	qsin_lut[0724] =  9'sd149;
	icos_lut[0724] =  9'sd149;
	qsin_lut[0725] =  9'sd175;
	icos_lut[0725] =  9'sd117;
	qsin_lut[0726] =  9'sd195;
	icos_lut[0726] =  9'sd81;
	qsin_lut[0727] =  9'sd207;
	icos_lut[0727] =  9'sd41;
	qsin_lut[0728] =  9'sd211;
	icos_lut[0728] =  9'sd0;
	qsin_lut[0729] =  9'sd207;
	icos_lut[0729] = -9'sd41;
	qsin_lut[0730] =  9'sd195;
	icos_lut[0730] = -9'sd81;
	qsin_lut[0731] =  9'sd175;
	icos_lut[0731] = -9'sd117;
	qsin_lut[0732] =  9'sd149;
	icos_lut[0732] = -9'sd149;
	qsin_lut[0733] =  9'sd117;
	icos_lut[0733] = -9'sd175;
	qsin_lut[0734] =  9'sd81;
	icos_lut[0734] = -9'sd195;
	qsin_lut[0735] =  9'sd41;
	icos_lut[0735] = -9'sd207;
	qsin_lut[0736] =  9'sd0;
	icos_lut[0736] = -9'sd209;
	qsin_lut[0737] = -9'sd41;
	icos_lut[0737] = -9'sd205;
	qsin_lut[0738] = -9'sd80;
	icos_lut[0738] = -9'sd193;
	qsin_lut[0739] = -9'sd116;
	icos_lut[0739] = -9'sd174;
	qsin_lut[0740] = -9'sd148;
	icos_lut[0740] = -9'sd148;
	qsin_lut[0741] = -9'sd174;
	icos_lut[0741] = -9'sd116;
	qsin_lut[0742] = -9'sd193;
	icos_lut[0742] = -9'sd80;
	qsin_lut[0743] = -9'sd205;
	icos_lut[0743] = -9'sd41;
	qsin_lut[0744] = -9'sd209;
	icos_lut[0744] = -9'sd0;
	qsin_lut[0745] = -9'sd205;
	icos_lut[0745] =  9'sd41;
	qsin_lut[0746] = -9'sd193;
	icos_lut[0746] =  9'sd80;
	qsin_lut[0747] = -9'sd174;
	icos_lut[0747] =  9'sd116;
	qsin_lut[0748] = -9'sd148;
	icos_lut[0748] =  9'sd148;
	qsin_lut[0749] = -9'sd116;
	icos_lut[0749] =  9'sd174;
	qsin_lut[0750] = -9'sd80;
	icos_lut[0750] =  9'sd193;
	qsin_lut[0751] = -9'sd41;
	icos_lut[0751] =  9'sd205;
	qsin_lut[0752] = -9'sd0;
	icos_lut[0752] =  9'sd209;
	qsin_lut[0753] =  9'sd41;
	icos_lut[0753] =  9'sd205;
	qsin_lut[0754] =  9'sd80;
	icos_lut[0754] =  9'sd193;
	qsin_lut[0755] =  9'sd116;
	icos_lut[0755] =  9'sd174;
	qsin_lut[0756] =  9'sd148;
	icos_lut[0756] =  9'sd148;
	qsin_lut[0757] =  9'sd174;
	icos_lut[0757] =  9'sd116;
	qsin_lut[0758] =  9'sd193;
	icos_lut[0758] =  9'sd80;
	qsin_lut[0759] =  9'sd205;
	icos_lut[0759] =  9'sd41;
	qsin_lut[0760] =  9'sd209;
	icos_lut[0760] =  9'sd0;
	qsin_lut[0761] =  9'sd205;
	icos_lut[0761] = -9'sd41;
	qsin_lut[0762] =  9'sd193;
	icos_lut[0762] = -9'sd80;
	qsin_lut[0763] =  9'sd174;
	icos_lut[0763] = -9'sd116;
	qsin_lut[0764] =  9'sd148;
	icos_lut[0764] = -9'sd148;
	qsin_lut[0765] =  9'sd116;
	icos_lut[0765] = -9'sd174;
	qsin_lut[0766] =  9'sd80;
	icos_lut[0766] = -9'sd193;
	qsin_lut[0767] =  9'sd41;
	icos_lut[0767] = -9'sd205;
	qsin_lut[0768] =  9'sd0;
	icos_lut[0768] = -9'sd207;
	qsin_lut[0769] = -9'sd40;
	icos_lut[0769] = -9'sd203;
	qsin_lut[0770] = -9'sd79;
	icos_lut[0770] = -9'sd191;
	qsin_lut[0771] = -9'sd115;
	icos_lut[0771] = -9'sd172;
	qsin_lut[0772] = -9'sd146;
	icos_lut[0772] = -9'sd146;
	qsin_lut[0773] = -9'sd172;
	icos_lut[0773] = -9'sd115;
	qsin_lut[0774] = -9'sd191;
	icos_lut[0774] = -9'sd79;
	qsin_lut[0775] = -9'sd203;
	icos_lut[0775] = -9'sd40;
	qsin_lut[0776] = -9'sd207;
	icos_lut[0776] = -9'sd0;
	qsin_lut[0777] = -9'sd203;
	icos_lut[0777] =  9'sd40;
	qsin_lut[0778] = -9'sd191;
	icos_lut[0778] =  9'sd79;
	qsin_lut[0779] = -9'sd172;
	icos_lut[0779] =  9'sd115;
	qsin_lut[0780] = -9'sd146;
	icos_lut[0780] =  9'sd146;
	qsin_lut[0781] = -9'sd115;
	icos_lut[0781] =  9'sd172;
	qsin_lut[0782] = -9'sd79;
	icos_lut[0782] =  9'sd191;
	qsin_lut[0783] = -9'sd40;
	icos_lut[0783] =  9'sd203;
	qsin_lut[0784] = -9'sd0;
	icos_lut[0784] =  9'sd207;
	qsin_lut[0785] =  9'sd40;
	icos_lut[0785] =  9'sd203;
	qsin_lut[0786] =  9'sd79;
	icos_lut[0786] =  9'sd191;
	qsin_lut[0787] =  9'sd115;
	icos_lut[0787] =  9'sd172;
	qsin_lut[0788] =  9'sd146;
	icos_lut[0788] =  9'sd146;
	qsin_lut[0789] =  9'sd172;
	icos_lut[0789] =  9'sd115;
	qsin_lut[0790] =  9'sd191;
	icos_lut[0790] =  9'sd79;
	qsin_lut[0791] =  9'sd203;
	icos_lut[0791] =  9'sd40;
	qsin_lut[0792] =  9'sd207;
	icos_lut[0792] =  9'sd0;
	qsin_lut[0793] =  9'sd203;
	icos_lut[0793] = -9'sd40;
	qsin_lut[0794] =  9'sd191;
	icos_lut[0794] = -9'sd79;
	qsin_lut[0795] =  9'sd172;
	icos_lut[0795] = -9'sd115;
	qsin_lut[0796] =  9'sd146;
	icos_lut[0796] = -9'sd146;
	qsin_lut[0797] =  9'sd115;
	icos_lut[0797] = -9'sd172;
	qsin_lut[0798] =  9'sd79;
	icos_lut[0798] = -9'sd191;
	qsin_lut[0799] =  9'sd40;
	icos_lut[0799] = -9'sd203;
	qsin_lut[0800] =  9'sd0;
	icos_lut[0800] = -9'sd205;
	qsin_lut[0801] = -9'sd40;
	icos_lut[0801] = -9'sd201;
	qsin_lut[0802] = -9'sd78;
	icos_lut[0802] = -9'sd189;
	qsin_lut[0803] = -9'sd114;
	icos_lut[0803] = -9'sd170;
	qsin_lut[0804] = -9'sd145;
	icos_lut[0804] = -9'sd145;
	qsin_lut[0805] = -9'sd170;
	icos_lut[0805] = -9'sd114;
	qsin_lut[0806] = -9'sd189;
	icos_lut[0806] = -9'sd78;
	qsin_lut[0807] = -9'sd201;
	icos_lut[0807] = -9'sd40;
	qsin_lut[0808] = -9'sd205;
	icos_lut[0808] = -9'sd0;
	qsin_lut[0809] = -9'sd201;
	icos_lut[0809] =  9'sd40;
	qsin_lut[0810] = -9'sd189;
	icos_lut[0810] =  9'sd78;
	qsin_lut[0811] = -9'sd170;
	icos_lut[0811] =  9'sd114;
	qsin_lut[0812] = -9'sd145;
	icos_lut[0812] =  9'sd145;
	qsin_lut[0813] = -9'sd114;
	icos_lut[0813] =  9'sd170;
	qsin_lut[0814] = -9'sd78;
	icos_lut[0814] =  9'sd189;
	qsin_lut[0815] = -9'sd40;
	icos_lut[0815] =  9'sd201;
	qsin_lut[0816] = -9'sd0;
	icos_lut[0816] =  9'sd205;
	qsin_lut[0817] =  9'sd40;
	icos_lut[0817] =  9'sd201;
	qsin_lut[0818] =  9'sd78;
	icos_lut[0818] =  9'sd189;
	qsin_lut[0819] =  9'sd114;
	icos_lut[0819] =  9'sd170;
	qsin_lut[0820] =  9'sd145;
	icos_lut[0820] =  9'sd145;
	qsin_lut[0821] =  9'sd170;
	icos_lut[0821] =  9'sd114;
	qsin_lut[0822] =  9'sd189;
	icos_lut[0822] =  9'sd78;
	qsin_lut[0823] =  9'sd201;
	icos_lut[0823] =  9'sd40;
	qsin_lut[0824] =  9'sd205;
	icos_lut[0824] =  9'sd0;
	qsin_lut[0825] =  9'sd201;
	icos_lut[0825] = -9'sd40;
	qsin_lut[0826] =  9'sd189;
	icos_lut[0826] = -9'sd78;
	qsin_lut[0827] =  9'sd170;
	icos_lut[0827] = -9'sd114;
	qsin_lut[0828] =  9'sd145;
	icos_lut[0828] = -9'sd145;
	qsin_lut[0829] =  9'sd114;
	icos_lut[0829] = -9'sd170;
	qsin_lut[0830] =  9'sd78;
	icos_lut[0830] = -9'sd189;
	qsin_lut[0831] =  9'sd40;
	icos_lut[0831] = -9'sd201;
	qsin_lut[0832] =  9'sd0;
	icos_lut[0832] = -9'sd203;
	qsin_lut[0833] = -9'sd40;
	icos_lut[0833] = -9'sd199;
	qsin_lut[0834] = -9'sd78;
	icos_lut[0834] = -9'sd188;
	qsin_lut[0835] = -9'sd113;
	icos_lut[0835] = -9'sd169;
	qsin_lut[0836] = -9'sd144;
	icos_lut[0836] = -9'sd144;
	qsin_lut[0837] = -9'sd169;
	icos_lut[0837] = -9'sd113;
	qsin_lut[0838] = -9'sd188;
	icos_lut[0838] = -9'sd78;
	qsin_lut[0839] = -9'sd199;
	icos_lut[0839] = -9'sd40;
	qsin_lut[0840] = -9'sd203;
	icos_lut[0840] = -9'sd0;
	qsin_lut[0841] = -9'sd199;
	icos_lut[0841] =  9'sd40;
	qsin_lut[0842] = -9'sd188;
	icos_lut[0842] =  9'sd78;
	qsin_lut[0843] = -9'sd169;
	icos_lut[0843] =  9'sd113;
	qsin_lut[0844] = -9'sd144;
	icos_lut[0844] =  9'sd144;
	qsin_lut[0845] = -9'sd113;
	icos_lut[0845] =  9'sd169;
	qsin_lut[0846] = -9'sd78;
	icos_lut[0846] =  9'sd188;
	qsin_lut[0847] = -9'sd40;
	icos_lut[0847] =  9'sd199;
	qsin_lut[0848] = -9'sd0;
	icos_lut[0848] =  9'sd203;
	qsin_lut[0849] =  9'sd40;
	icos_lut[0849] =  9'sd199;
	qsin_lut[0850] =  9'sd78;
	icos_lut[0850] =  9'sd188;
	qsin_lut[0851] =  9'sd113;
	icos_lut[0851] =  9'sd169;
	qsin_lut[0852] =  9'sd144;
	icos_lut[0852] =  9'sd144;
	qsin_lut[0853] =  9'sd169;
	icos_lut[0853] =  9'sd113;
	qsin_lut[0854] =  9'sd188;
	icos_lut[0854] =  9'sd78;
	qsin_lut[0855] =  9'sd199;
	icos_lut[0855] =  9'sd40;
	qsin_lut[0856] =  9'sd203;
	icos_lut[0856] =  9'sd0;
	qsin_lut[0857] =  9'sd199;
	icos_lut[0857] = -9'sd40;
	qsin_lut[0858] =  9'sd188;
	icos_lut[0858] = -9'sd78;
	qsin_lut[0859] =  9'sd169;
	icos_lut[0859] = -9'sd113;
	qsin_lut[0860] =  9'sd144;
	icos_lut[0860] = -9'sd144;
	qsin_lut[0861] =  9'sd113;
	icos_lut[0861] = -9'sd169;
	qsin_lut[0862] =  9'sd78;
	icos_lut[0862] = -9'sd188;
	qsin_lut[0863] =  9'sd40;
	icos_lut[0863] = -9'sd199;
	qsin_lut[0864] =  9'sd0;
	icos_lut[0864] = -9'sd201;
	qsin_lut[0865] = -9'sd39;
	icos_lut[0865] = -9'sd197;
	qsin_lut[0866] = -9'sd77;
	icos_lut[0866] = -9'sd186;
	qsin_lut[0867] = -9'sd112;
	icos_lut[0867] = -9'sd167;
	qsin_lut[0868] = -9'sd142;
	icos_lut[0868] = -9'sd142;
	qsin_lut[0869] = -9'sd167;
	icos_lut[0869] = -9'sd112;
	qsin_lut[0870] = -9'sd186;
	icos_lut[0870] = -9'sd77;
	qsin_lut[0871] = -9'sd197;
	icos_lut[0871] = -9'sd39;
	qsin_lut[0872] = -9'sd201;
	icos_lut[0872] = -9'sd0;
	qsin_lut[0873] = -9'sd197;
	icos_lut[0873] =  9'sd39;
	qsin_lut[0874] = -9'sd186;
	icos_lut[0874] =  9'sd77;
	qsin_lut[0875] = -9'sd167;
	icos_lut[0875] =  9'sd112;
	qsin_lut[0876] = -9'sd142;
	icos_lut[0876] =  9'sd142;
	qsin_lut[0877] = -9'sd112;
	icos_lut[0877] =  9'sd167;
	qsin_lut[0878] = -9'sd77;
	icos_lut[0878] =  9'sd186;
	qsin_lut[0879] = -9'sd39;
	icos_lut[0879] =  9'sd197;
	qsin_lut[0880] = -9'sd0;
	icos_lut[0880] =  9'sd201;
	qsin_lut[0881] =  9'sd39;
	icos_lut[0881] =  9'sd197;
	qsin_lut[0882] =  9'sd77;
	icos_lut[0882] =  9'sd186;
	qsin_lut[0883] =  9'sd112;
	icos_lut[0883] =  9'sd167;
	qsin_lut[0884] =  9'sd142;
	icos_lut[0884] =  9'sd142;
	qsin_lut[0885] =  9'sd167;
	icos_lut[0885] =  9'sd112;
	qsin_lut[0886] =  9'sd186;
	icos_lut[0886] =  9'sd77;
	qsin_lut[0887] =  9'sd197;
	icos_lut[0887] =  9'sd39;
	qsin_lut[0888] =  9'sd201;
	icos_lut[0888] =  9'sd0;
	qsin_lut[0889] =  9'sd197;
	icos_lut[0889] = -9'sd39;
	qsin_lut[0890] =  9'sd186;
	icos_lut[0890] = -9'sd77;
	qsin_lut[0891] =  9'sd167;
	icos_lut[0891] = -9'sd112;
	qsin_lut[0892] =  9'sd142;
	icos_lut[0892] = -9'sd142;
	qsin_lut[0893] =  9'sd112;
	icos_lut[0893] = -9'sd167;
	qsin_lut[0894] =  9'sd77;
	icos_lut[0894] = -9'sd186;
	qsin_lut[0895] =  9'sd39;
	icos_lut[0895] = -9'sd197;
	qsin_lut[0896] =  9'sd0;
	icos_lut[0896] = -9'sd199;
	qsin_lut[0897] = -9'sd39;
	icos_lut[0897] = -9'sd195;
	qsin_lut[0898] = -9'sd76;
	icos_lut[0898] = -9'sd184;
	qsin_lut[0899] = -9'sd111;
	icos_lut[0899] = -9'sd165;
	qsin_lut[0900] = -9'sd141;
	icos_lut[0900] = -9'sd141;
	qsin_lut[0901] = -9'sd165;
	icos_lut[0901] = -9'sd111;
	qsin_lut[0902] = -9'sd184;
	icos_lut[0902] = -9'sd76;
	qsin_lut[0903] = -9'sd195;
	icos_lut[0903] = -9'sd39;
	qsin_lut[0904] = -9'sd199;
	icos_lut[0904] = -9'sd0;
	qsin_lut[0905] = -9'sd195;
	icos_lut[0905] =  9'sd39;
	qsin_lut[0906] = -9'sd184;
	icos_lut[0906] =  9'sd76;
	qsin_lut[0907] = -9'sd165;
	icos_lut[0907] =  9'sd111;
	qsin_lut[0908] = -9'sd141;
	icos_lut[0908] =  9'sd141;
	qsin_lut[0909] = -9'sd111;
	icos_lut[0909] =  9'sd165;
	qsin_lut[0910] = -9'sd76;
	icos_lut[0910] =  9'sd184;
	qsin_lut[0911] = -9'sd39;
	icos_lut[0911] =  9'sd195;
	qsin_lut[0912] = -9'sd0;
	icos_lut[0912] =  9'sd199;
	qsin_lut[0913] =  9'sd39;
	icos_lut[0913] =  9'sd195;
	qsin_lut[0914] =  9'sd76;
	icos_lut[0914] =  9'sd184;
	qsin_lut[0915] =  9'sd111;
	icos_lut[0915] =  9'sd165;
	qsin_lut[0916] =  9'sd141;
	icos_lut[0916] =  9'sd141;
	qsin_lut[0917] =  9'sd165;
	icos_lut[0917] =  9'sd111;
	qsin_lut[0918] =  9'sd184;
	icos_lut[0918] =  9'sd76;
	qsin_lut[0919] =  9'sd195;
	icos_lut[0919] =  9'sd39;
	qsin_lut[0920] =  9'sd199;
	icos_lut[0920] =  9'sd0;
	qsin_lut[0921] =  9'sd195;
	icos_lut[0921] = -9'sd39;
	qsin_lut[0922] =  9'sd184;
	icos_lut[0922] = -9'sd76;
	qsin_lut[0923] =  9'sd165;
	icos_lut[0923] = -9'sd111;
	qsin_lut[0924] =  9'sd141;
	icos_lut[0924] = -9'sd141;
	qsin_lut[0925] =  9'sd111;
	icos_lut[0925] = -9'sd165;
	qsin_lut[0926] =  9'sd76;
	icos_lut[0926] = -9'sd184;
	qsin_lut[0927] =  9'sd39;
	icos_lut[0927] = -9'sd195;
	qsin_lut[0928] =  9'sd0;
	icos_lut[0928] = -9'sd197;
	qsin_lut[0929] = -9'sd38;
	icos_lut[0929] = -9'sd193;
	qsin_lut[0930] = -9'sd75;
	icos_lut[0930] = -9'sd182;
	qsin_lut[0931] = -9'sd109;
	icos_lut[0931] = -9'sd164;
	qsin_lut[0932] = -9'sd139;
	icos_lut[0932] = -9'sd139;
	qsin_lut[0933] = -9'sd164;
	icos_lut[0933] = -9'sd109;
	qsin_lut[0934] = -9'sd182;
	icos_lut[0934] = -9'sd75;
	qsin_lut[0935] = -9'sd193;
	icos_lut[0935] = -9'sd38;
	qsin_lut[0936] = -9'sd197;
	icos_lut[0936] = -9'sd0;
	qsin_lut[0937] = -9'sd193;
	icos_lut[0937] =  9'sd38;
	qsin_lut[0938] = -9'sd182;
	icos_lut[0938] =  9'sd75;
	qsin_lut[0939] = -9'sd164;
	icos_lut[0939] =  9'sd109;
	qsin_lut[0940] = -9'sd139;
	icos_lut[0940] =  9'sd139;
	qsin_lut[0941] = -9'sd109;
	icos_lut[0941] =  9'sd164;
	qsin_lut[0942] = -9'sd75;
	icos_lut[0942] =  9'sd182;
	qsin_lut[0943] = -9'sd38;
	icos_lut[0943] =  9'sd193;
	qsin_lut[0944] = -9'sd0;
	icos_lut[0944] =  9'sd197;
	qsin_lut[0945] =  9'sd38;
	icos_lut[0945] =  9'sd193;
	qsin_lut[0946] =  9'sd75;
	icos_lut[0946] =  9'sd182;
	qsin_lut[0947] =  9'sd109;
	icos_lut[0947] =  9'sd164;
	qsin_lut[0948] =  9'sd139;
	icos_lut[0948] =  9'sd139;
	qsin_lut[0949] =  9'sd164;
	icos_lut[0949] =  9'sd109;
	qsin_lut[0950] =  9'sd182;
	icos_lut[0950] =  9'sd75;
	qsin_lut[0951] =  9'sd193;
	icos_lut[0951] =  9'sd38;
	qsin_lut[0952] =  9'sd197;
	icos_lut[0952] =  9'sd0;
	qsin_lut[0953] =  9'sd193;
	icos_lut[0953] = -9'sd38;
	qsin_lut[0954] =  9'sd182;
	icos_lut[0954] = -9'sd75;
	qsin_lut[0955] =  9'sd164;
	icos_lut[0955] = -9'sd109;
	qsin_lut[0956] =  9'sd139;
	icos_lut[0956] = -9'sd139;
	qsin_lut[0957] =  9'sd109;
	icos_lut[0957] = -9'sd164;
	qsin_lut[0958] =  9'sd75;
	icos_lut[0958] = -9'sd182;
	qsin_lut[0959] =  9'sd38;
	icos_lut[0959] = -9'sd193;
	qsin_lut[0960] =  9'sd0;
	icos_lut[0960] = -9'sd195;
	qsin_lut[0961] = -9'sd38;
	icos_lut[0961] = -9'sd191;
	qsin_lut[0962] = -9'sd75;
	icos_lut[0962] = -9'sd180;
	qsin_lut[0963] = -9'sd108;
	icos_lut[0963] = -9'sd162;
	qsin_lut[0964] = -9'sd138;
	icos_lut[0964] = -9'sd138;
	qsin_lut[0965] = -9'sd162;
	icos_lut[0965] = -9'sd108;
	qsin_lut[0966] = -9'sd180;
	icos_lut[0966] = -9'sd75;
	qsin_lut[0967] = -9'sd191;
	icos_lut[0967] = -9'sd38;
	qsin_lut[0968] = -9'sd195;
	icos_lut[0968] = -9'sd0;
	qsin_lut[0969] = -9'sd191;
	icos_lut[0969] =  9'sd38;
	qsin_lut[0970] = -9'sd180;
	icos_lut[0970] =  9'sd75;
	qsin_lut[0971] = -9'sd162;
	icos_lut[0971] =  9'sd108;
	qsin_lut[0972] = -9'sd138;
	icos_lut[0972] =  9'sd138;
	qsin_lut[0973] = -9'sd108;
	icos_lut[0973] =  9'sd162;
	qsin_lut[0974] = -9'sd75;
	icos_lut[0974] =  9'sd180;
	qsin_lut[0975] = -9'sd38;
	icos_lut[0975] =  9'sd191;
	qsin_lut[0976] = -9'sd0;
	icos_lut[0976] =  9'sd195;
	qsin_lut[0977] =  9'sd38;
	icos_lut[0977] =  9'sd191;
	qsin_lut[0978] =  9'sd75;
	icos_lut[0978] =  9'sd180;
	qsin_lut[0979] =  9'sd108;
	icos_lut[0979] =  9'sd162;
	qsin_lut[0980] =  9'sd138;
	icos_lut[0980] =  9'sd138;
	qsin_lut[0981] =  9'sd162;
	icos_lut[0981] =  9'sd108;
	qsin_lut[0982] =  9'sd180;
	icos_lut[0982] =  9'sd75;
	qsin_lut[0983] =  9'sd191;
	icos_lut[0983] =  9'sd38;
	qsin_lut[0984] =  9'sd195;
	icos_lut[0984] =  9'sd0;
	qsin_lut[0985] =  9'sd191;
	icos_lut[0985] = -9'sd38;
	qsin_lut[0986] =  9'sd180;
	icos_lut[0986] = -9'sd75;
	qsin_lut[0987] =  9'sd162;
	icos_lut[0987] = -9'sd108;
	qsin_lut[0988] =  9'sd138;
	icos_lut[0988] = -9'sd138;
	qsin_lut[0989] =  9'sd108;
	icos_lut[0989] = -9'sd162;
	qsin_lut[0990] =  9'sd75;
	icos_lut[0990] = -9'sd180;
	qsin_lut[0991] =  9'sd38;
	icos_lut[0991] = -9'sd191;
	qsin_lut[0992] =  9'sd0;
	icos_lut[0992] = -9'sd193;
	qsin_lut[0993] = -9'sd38;
	icos_lut[0993] = -9'sd189;
	qsin_lut[0994] = -9'sd74;
	icos_lut[0994] = -9'sd178;
	qsin_lut[0995] = -9'sd107;
	icos_lut[0995] = -9'sd160;
	qsin_lut[0996] = -9'sd136;
	icos_lut[0996] = -9'sd136;
	qsin_lut[0997] = -9'sd160;
	icos_lut[0997] = -9'sd107;
	qsin_lut[0998] = -9'sd178;
	icos_lut[0998] = -9'sd74;
	qsin_lut[0999] = -9'sd189;
	icos_lut[0999] = -9'sd38;
	qsin_lut[1000] = -9'sd193;
	icos_lut[1000] = -9'sd0;
	qsin_lut[1001] = -9'sd189;
	icos_lut[1001] =  9'sd38;
	qsin_lut[1002] = -9'sd178;
	icos_lut[1002] =  9'sd74;
	qsin_lut[1003] = -9'sd160;
	icos_lut[1003] =  9'sd107;
	qsin_lut[1004] = -9'sd136;
	icos_lut[1004] =  9'sd136;
	qsin_lut[1005] = -9'sd107;
	icos_lut[1005] =  9'sd160;
	qsin_lut[1006] = -9'sd74;
	icos_lut[1006] =  9'sd178;
	qsin_lut[1007] = -9'sd38;
	icos_lut[1007] =  9'sd189;
	qsin_lut[1008] = -9'sd0;
	icos_lut[1008] =  9'sd193;
	qsin_lut[1009] =  9'sd38;
	icos_lut[1009] =  9'sd189;
	qsin_lut[1010] =  9'sd74;
	icos_lut[1010] =  9'sd178;
	qsin_lut[1011] =  9'sd107;
	icos_lut[1011] =  9'sd160;
	qsin_lut[1012] =  9'sd136;
	icos_lut[1012] =  9'sd136;
	qsin_lut[1013] =  9'sd160;
	icos_lut[1013] =  9'sd107;
	qsin_lut[1014] =  9'sd178;
	icos_lut[1014] =  9'sd74;
	qsin_lut[1015] =  9'sd189;
	icos_lut[1015] =  9'sd38;
	qsin_lut[1016] =  9'sd193;
	icos_lut[1016] =  9'sd0;
	qsin_lut[1017] =  9'sd189;
	icos_lut[1017] = -9'sd38;
	qsin_lut[1018] =  9'sd178;
	icos_lut[1018] = -9'sd74;
	qsin_lut[1019] =  9'sd160;
	icos_lut[1019] = -9'sd107;
	qsin_lut[1020] =  9'sd136;
	icos_lut[1020] = -9'sd136;
	qsin_lut[1021] =  9'sd107;
	icos_lut[1021] = -9'sd160;
	qsin_lut[1022] =  9'sd74;
	icos_lut[1022] = -9'sd178;
	qsin_lut[1023] =  9'sd38;
	icos_lut[1023] = -9'sd189;
	qsin_lut[1024] =  9'sd0;
	icos_lut[1024] = -9'sd191;
	qsin_lut[1025] = -9'sd37;
	icos_lut[1025] = -9'sd187;
	qsin_lut[1026] = -9'sd73;
	icos_lut[1026] = -9'sd176;
	qsin_lut[1027] = -9'sd106;
	icos_lut[1027] = -9'sd159;
	qsin_lut[1028] = -9'sd135;
	icos_lut[1028] = -9'sd135;
	qsin_lut[1029] = -9'sd159;
	icos_lut[1029] = -9'sd106;
	qsin_lut[1030] = -9'sd176;
	icos_lut[1030] = -9'sd73;
	qsin_lut[1031] = -9'sd187;
	icos_lut[1031] = -9'sd37;
	qsin_lut[1032] = -9'sd191;
	icos_lut[1032] = -9'sd0;
	qsin_lut[1033] = -9'sd187;
	icos_lut[1033] =  9'sd37;
	qsin_lut[1034] = -9'sd176;
	icos_lut[1034] =  9'sd73;
	qsin_lut[1035] = -9'sd159;
	icos_lut[1035] =  9'sd106;
	qsin_lut[1036] = -9'sd135;
	icos_lut[1036] =  9'sd135;
	qsin_lut[1037] = -9'sd106;
	icos_lut[1037] =  9'sd159;
	qsin_lut[1038] = -9'sd73;
	icos_lut[1038] =  9'sd176;
	qsin_lut[1039] = -9'sd37;
	icos_lut[1039] =  9'sd187;
	qsin_lut[1040] = -9'sd0;
	icos_lut[1040] =  9'sd191;
	qsin_lut[1041] =  9'sd37;
	icos_lut[1041] =  9'sd187;
	qsin_lut[1042] =  9'sd73;
	icos_lut[1042] =  9'sd176;
	qsin_lut[1043] =  9'sd106;
	icos_lut[1043] =  9'sd159;
	qsin_lut[1044] =  9'sd135;
	icos_lut[1044] =  9'sd135;
	qsin_lut[1045] =  9'sd159;
	icos_lut[1045] =  9'sd106;
	qsin_lut[1046] =  9'sd176;
	icos_lut[1046] =  9'sd73;
	qsin_lut[1047] =  9'sd187;
	icos_lut[1047] =  9'sd37;
	qsin_lut[1048] =  9'sd191;
	icos_lut[1048] =  9'sd0;
	qsin_lut[1049] =  9'sd187;
	icos_lut[1049] = -9'sd37;
	qsin_lut[1050] =  9'sd176;
	icos_lut[1050] = -9'sd73;
	qsin_lut[1051] =  9'sd159;
	icos_lut[1051] = -9'sd106;
	qsin_lut[1052] =  9'sd135;
	icos_lut[1052] = -9'sd135;
	qsin_lut[1053] =  9'sd106;
	icos_lut[1053] = -9'sd159;
	qsin_lut[1054] =  9'sd73;
	icos_lut[1054] = -9'sd176;
	qsin_lut[1055] =  9'sd37;
	icos_lut[1055] = -9'sd187;
	qsin_lut[1056] =  9'sd0;
	icos_lut[1056] = -9'sd189;
	qsin_lut[1057] = -9'sd37;
	icos_lut[1057] = -9'sd185;
	qsin_lut[1058] = -9'sd72;
	icos_lut[1058] = -9'sd175;
	qsin_lut[1059] = -9'sd105;
	icos_lut[1059] = -9'sd157;
	qsin_lut[1060] = -9'sd134;
	icos_lut[1060] = -9'sd134;
	qsin_lut[1061] = -9'sd157;
	icos_lut[1061] = -9'sd105;
	qsin_lut[1062] = -9'sd175;
	icos_lut[1062] = -9'sd72;
	qsin_lut[1063] = -9'sd185;
	icos_lut[1063] = -9'sd37;
	qsin_lut[1064] = -9'sd189;
	icos_lut[1064] = -9'sd0;
	qsin_lut[1065] = -9'sd185;
	icos_lut[1065] =  9'sd37;
	qsin_lut[1066] = -9'sd175;
	icos_lut[1066] =  9'sd72;
	qsin_lut[1067] = -9'sd157;
	icos_lut[1067] =  9'sd105;
	qsin_lut[1068] = -9'sd134;
	icos_lut[1068] =  9'sd134;
	qsin_lut[1069] = -9'sd105;
	icos_lut[1069] =  9'sd157;
	qsin_lut[1070] = -9'sd72;
	icos_lut[1070] =  9'sd175;
	qsin_lut[1071] = -9'sd37;
	icos_lut[1071] =  9'sd185;
	qsin_lut[1072] = -9'sd0;
	icos_lut[1072] =  9'sd189;
	qsin_lut[1073] =  9'sd37;
	icos_lut[1073] =  9'sd185;
	qsin_lut[1074] =  9'sd72;
	icos_lut[1074] =  9'sd175;
	qsin_lut[1075] =  9'sd105;
	icos_lut[1075] =  9'sd157;
	qsin_lut[1076] =  9'sd134;
	icos_lut[1076] =  9'sd134;
	qsin_lut[1077] =  9'sd157;
	icos_lut[1077] =  9'sd105;
	qsin_lut[1078] =  9'sd175;
	icos_lut[1078] =  9'sd72;
	qsin_lut[1079] =  9'sd185;
	icos_lut[1079] =  9'sd37;
	qsin_lut[1080] =  9'sd189;
	icos_lut[1080] =  9'sd0;
	qsin_lut[1081] =  9'sd185;
	icos_lut[1081] = -9'sd37;
	qsin_lut[1082] =  9'sd175;
	icos_lut[1082] = -9'sd72;
	qsin_lut[1083] =  9'sd157;
	icos_lut[1083] = -9'sd105;
	qsin_lut[1084] =  9'sd134;
	icos_lut[1084] = -9'sd134;
	qsin_lut[1085] =  9'sd105;
	icos_lut[1085] = -9'sd157;
	qsin_lut[1086] =  9'sd72;
	icos_lut[1086] = -9'sd175;
	qsin_lut[1087] =  9'sd37;
	icos_lut[1087] = -9'sd185;
	qsin_lut[1088] =  9'sd0;
	icos_lut[1088] = -9'sd187;
	qsin_lut[1089] = -9'sd36;
	icos_lut[1089] = -9'sd183;
	qsin_lut[1090] = -9'sd72;
	icos_lut[1090] = -9'sd173;
	qsin_lut[1091] = -9'sd104;
	icos_lut[1091] = -9'sd155;
	qsin_lut[1092] = -9'sd132;
	icos_lut[1092] = -9'sd132;
	qsin_lut[1093] = -9'sd155;
	icos_lut[1093] = -9'sd104;
	qsin_lut[1094] = -9'sd173;
	icos_lut[1094] = -9'sd72;
	qsin_lut[1095] = -9'sd183;
	icos_lut[1095] = -9'sd36;
	qsin_lut[1096] = -9'sd187;
	icos_lut[1096] = -9'sd0;
	qsin_lut[1097] = -9'sd183;
	icos_lut[1097] =  9'sd36;
	qsin_lut[1098] = -9'sd173;
	icos_lut[1098] =  9'sd72;
	qsin_lut[1099] = -9'sd155;
	icos_lut[1099] =  9'sd104;
	qsin_lut[1100] = -9'sd132;
	icos_lut[1100] =  9'sd132;
	qsin_lut[1101] = -9'sd104;
	icos_lut[1101] =  9'sd155;
	qsin_lut[1102] = -9'sd72;
	icos_lut[1102] =  9'sd173;
	qsin_lut[1103] = -9'sd36;
	icos_lut[1103] =  9'sd183;
	qsin_lut[1104] = -9'sd0;
	icos_lut[1104] =  9'sd187;
	qsin_lut[1105] =  9'sd36;
	icos_lut[1105] =  9'sd183;
	qsin_lut[1106] =  9'sd72;
	icos_lut[1106] =  9'sd173;
	qsin_lut[1107] =  9'sd104;
	icos_lut[1107] =  9'sd155;
	qsin_lut[1108] =  9'sd132;
	icos_lut[1108] =  9'sd132;
	qsin_lut[1109] =  9'sd155;
	icos_lut[1109] =  9'sd104;
	qsin_lut[1110] =  9'sd173;
	icos_lut[1110] =  9'sd72;
	qsin_lut[1111] =  9'sd183;
	icos_lut[1111] =  9'sd36;
	qsin_lut[1112] =  9'sd187;
	icos_lut[1112] =  9'sd0;
	qsin_lut[1113] =  9'sd183;
	icos_lut[1113] = -9'sd36;
	qsin_lut[1114] =  9'sd173;
	icos_lut[1114] = -9'sd72;
	qsin_lut[1115] =  9'sd155;
	icos_lut[1115] = -9'sd104;
	qsin_lut[1116] =  9'sd132;
	icos_lut[1116] = -9'sd132;
	qsin_lut[1117] =  9'sd104;
	icos_lut[1117] = -9'sd155;
	qsin_lut[1118] =  9'sd72;
	icos_lut[1118] = -9'sd173;
	qsin_lut[1119] =  9'sd36;
	icos_lut[1119] = -9'sd183;
	qsin_lut[1120] =  9'sd0;
	icos_lut[1120] = -9'sd185;
	qsin_lut[1121] = -9'sd36;
	icos_lut[1121] = -9'sd181;
	qsin_lut[1122] = -9'sd71;
	icos_lut[1122] = -9'sd171;
	qsin_lut[1123] = -9'sd103;
	icos_lut[1123] = -9'sd154;
	qsin_lut[1124] = -9'sd131;
	icos_lut[1124] = -9'sd131;
	qsin_lut[1125] = -9'sd154;
	icos_lut[1125] = -9'sd103;
	qsin_lut[1126] = -9'sd171;
	icos_lut[1126] = -9'sd71;
	qsin_lut[1127] = -9'sd181;
	icos_lut[1127] = -9'sd36;
	qsin_lut[1128] = -9'sd185;
	icos_lut[1128] = -9'sd0;
	qsin_lut[1129] = -9'sd181;
	icos_lut[1129] =  9'sd36;
	qsin_lut[1130] = -9'sd171;
	icos_lut[1130] =  9'sd71;
	qsin_lut[1131] = -9'sd154;
	icos_lut[1131] =  9'sd103;
	qsin_lut[1132] = -9'sd131;
	icos_lut[1132] =  9'sd131;
	qsin_lut[1133] = -9'sd103;
	icos_lut[1133] =  9'sd154;
	qsin_lut[1134] = -9'sd71;
	icos_lut[1134] =  9'sd171;
	qsin_lut[1135] = -9'sd36;
	icos_lut[1135] =  9'sd181;
	qsin_lut[1136] = -9'sd0;
	icos_lut[1136] =  9'sd185;
	qsin_lut[1137] =  9'sd36;
	icos_lut[1137] =  9'sd181;
	qsin_lut[1138] =  9'sd71;
	icos_lut[1138] =  9'sd171;
	qsin_lut[1139] =  9'sd103;
	icos_lut[1139] =  9'sd154;
	qsin_lut[1140] =  9'sd131;
	icos_lut[1140] =  9'sd131;
	qsin_lut[1141] =  9'sd154;
	icos_lut[1141] =  9'sd103;
	qsin_lut[1142] =  9'sd171;
	icos_lut[1142] =  9'sd71;
	qsin_lut[1143] =  9'sd181;
	icos_lut[1143] =  9'sd36;
	qsin_lut[1144] =  9'sd185;
	icos_lut[1144] =  9'sd0;
	qsin_lut[1145] =  9'sd181;
	icos_lut[1145] = -9'sd36;
	qsin_lut[1146] =  9'sd171;
	icos_lut[1146] = -9'sd71;
	qsin_lut[1147] =  9'sd154;
	icos_lut[1147] = -9'sd103;
	qsin_lut[1148] =  9'sd131;
	icos_lut[1148] = -9'sd131;
	qsin_lut[1149] =  9'sd103;
	icos_lut[1149] = -9'sd154;
	qsin_lut[1150] =  9'sd71;
	icos_lut[1150] = -9'sd171;
	qsin_lut[1151] =  9'sd36;
	icos_lut[1151] = -9'sd181;
	qsin_lut[1152] =  9'sd0;
	icos_lut[1152] = -9'sd183;
	qsin_lut[1153] = -9'sd36;
	icos_lut[1153] = -9'sd179;
	qsin_lut[1154] = -9'sd70;
	icos_lut[1154] = -9'sd169;
	qsin_lut[1155] = -9'sd102;
	icos_lut[1155] = -9'sd152;
	qsin_lut[1156] = -9'sd129;
	icos_lut[1156] = -9'sd129;
	qsin_lut[1157] = -9'sd152;
	icos_lut[1157] = -9'sd102;
	qsin_lut[1158] = -9'sd169;
	icos_lut[1158] = -9'sd70;
	qsin_lut[1159] = -9'sd179;
	icos_lut[1159] = -9'sd36;
	qsin_lut[1160] = -9'sd183;
	icos_lut[1160] = -9'sd0;
	qsin_lut[1161] = -9'sd179;
	icos_lut[1161] =  9'sd36;
	qsin_lut[1162] = -9'sd169;
	icos_lut[1162] =  9'sd70;
	qsin_lut[1163] = -9'sd152;
	icos_lut[1163] =  9'sd102;
	qsin_lut[1164] = -9'sd129;
	icos_lut[1164] =  9'sd129;
	qsin_lut[1165] = -9'sd102;
	icos_lut[1165] =  9'sd152;
	qsin_lut[1166] = -9'sd70;
	icos_lut[1166] =  9'sd169;
	qsin_lut[1167] = -9'sd36;
	icos_lut[1167] =  9'sd179;
	qsin_lut[1168] = -9'sd0;
	icos_lut[1168] =  9'sd183;
	qsin_lut[1169] =  9'sd36;
	icos_lut[1169] =  9'sd179;
	qsin_lut[1170] =  9'sd70;
	icos_lut[1170] =  9'sd169;
	qsin_lut[1171] =  9'sd102;
	icos_lut[1171] =  9'sd152;
	qsin_lut[1172] =  9'sd129;
	icos_lut[1172] =  9'sd129;
	qsin_lut[1173] =  9'sd152;
	icos_lut[1173] =  9'sd102;
	qsin_lut[1174] =  9'sd169;
	icos_lut[1174] =  9'sd70;
	qsin_lut[1175] =  9'sd179;
	icos_lut[1175] =  9'sd36;
	qsin_lut[1176] =  9'sd183;
	icos_lut[1176] =  9'sd0;
	qsin_lut[1177] =  9'sd179;
	icos_lut[1177] = -9'sd36;
	qsin_lut[1178] =  9'sd169;
	icos_lut[1178] = -9'sd70;
	qsin_lut[1179] =  9'sd152;
	icos_lut[1179] = -9'sd102;
	qsin_lut[1180] =  9'sd129;
	icos_lut[1180] = -9'sd129;
	qsin_lut[1181] =  9'sd102;
	icos_lut[1181] = -9'sd152;
	qsin_lut[1182] =  9'sd70;
	icos_lut[1182] = -9'sd169;
	qsin_lut[1183] =  9'sd36;
	icos_lut[1183] = -9'sd179;
	qsin_lut[1184] =  9'sd0;
	icos_lut[1184] = -9'sd181;
	qsin_lut[1185] = -9'sd35;
	icos_lut[1185] = -9'sd178;
	qsin_lut[1186] = -9'sd69;
	icos_lut[1186] = -9'sd167;
	qsin_lut[1187] = -9'sd101;
	icos_lut[1187] = -9'sd150;
	qsin_lut[1188] = -9'sd128;
	icos_lut[1188] = -9'sd128;
	qsin_lut[1189] = -9'sd150;
	icos_lut[1189] = -9'sd101;
	qsin_lut[1190] = -9'sd167;
	icos_lut[1190] = -9'sd69;
	qsin_lut[1191] = -9'sd178;
	icos_lut[1191] = -9'sd35;
	qsin_lut[1192] = -9'sd181;
	icos_lut[1192] = -9'sd0;
	qsin_lut[1193] = -9'sd178;
	icos_lut[1193] =  9'sd35;
	qsin_lut[1194] = -9'sd167;
	icos_lut[1194] =  9'sd69;
	qsin_lut[1195] = -9'sd150;
	icos_lut[1195] =  9'sd101;
	qsin_lut[1196] = -9'sd128;
	icos_lut[1196] =  9'sd128;
	qsin_lut[1197] = -9'sd101;
	icos_lut[1197] =  9'sd150;
	qsin_lut[1198] = -9'sd69;
	icos_lut[1198] =  9'sd167;
	qsin_lut[1199] = -9'sd35;
	icos_lut[1199] =  9'sd178;
	qsin_lut[1200] = -9'sd0;
	icos_lut[1200] =  9'sd181;
	qsin_lut[1201] =  9'sd35;
	icos_lut[1201] =  9'sd178;
	qsin_lut[1202] =  9'sd69;
	icos_lut[1202] =  9'sd167;
	qsin_lut[1203] =  9'sd101;
	icos_lut[1203] =  9'sd150;
	qsin_lut[1204] =  9'sd128;
	icos_lut[1204] =  9'sd128;
	qsin_lut[1205] =  9'sd150;
	icos_lut[1205] =  9'sd101;
	qsin_lut[1206] =  9'sd167;
	icos_lut[1206] =  9'sd69;
	qsin_lut[1207] =  9'sd178;
	icos_lut[1207] =  9'sd35;
	qsin_lut[1208] =  9'sd181;
	icos_lut[1208] =  9'sd0;
	qsin_lut[1209] =  9'sd178;
	icos_lut[1209] = -9'sd35;
	qsin_lut[1210] =  9'sd167;
	icos_lut[1210] = -9'sd69;
	qsin_lut[1211] =  9'sd150;
	icos_lut[1211] = -9'sd101;
	qsin_lut[1212] =  9'sd128;
	icos_lut[1212] = -9'sd128;
	qsin_lut[1213] =  9'sd101;
	icos_lut[1213] = -9'sd150;
	qsin_lut[1214] =  9'sd69;
	icos_lut[1214] = -9'sd167;
	qsin_lut[1215] =  9'sd35;
	icos_lut[1215] = -9'sd178;
	qsin_lut[1216] =  9'sd0;
	icos_lut[1216] = -9'sd179;
	qsin_lut[1217] = -9'sd35;
	icos_lut[1217] = -9'sd176;
	qsin_lut[1218] = -9'sd69;
	icos_lut[1218] = -9'sd165;
	qsin_lut[1219] = -9'sd99;
	icos_lut[1219] = -9'sd149;
	qsin_lut[1220] = -9'sd127;
	icos_lut[1220] = -9'sd127;
	qsin_lut[1221] = -9'sd149;
	icos_lut[1221] = -9'sd99;
	qsin_lut[1222] = -9'sd165;
	icos_lut[1222] = -9'sd69;
	qsin_lut[1223] = -9'sd176;
	icos_lut[1223] = -9'sd35;
	qsin_lut[1224] = -9'sd179;
	icos_lut[1224] = -9'sd0;
	qsin_lut[1225] = -9'sd176;
	icos_lut[1225] =  9'sd35;
	qsin_lut[1226] = -9'sd165;
	icos_lut[1226] =  9'sd69;
	qsin_lut[1227] = -9'sd149;
	icos_lut[1227] =  9'sd99;
	qsin_lut[1228] = -9'sd127;
	icos_lut[1228] =  9'sd127;
	qsin_lut[1229] = -9'sd99;
	icos_lut[1229] =  9'sd149;
	qsin_lut[1230] = -9'sd69;
	icos_lut[1230] =  9'sd165;
	qsin_lut[1231] = -9'sd35;
	icos_lut[1231] =  9'sd176;
	qsin_lut[1232] = -9'sd0;
	icos_lut[1232] =  9'sd179;
	qsin_lut[1233] =  9'sd35;
	icos_lut[1233] =  9'sd176;
	qsin_lut[1234] =  9'sd69;
	icos_lut[1234] =  9'sd165;
	qsin_lut[1235] =  9'sd99;
	icos_lut[1235] =  9'sd149;
	qsin_lut[1236] =  9'sd127;
	icos_lut[1236] =  9'sd127;
	qsin_lut[1237] =  9'sd149;
	icos_lut[1237] =  9'sd99;
	qsin_lut[1238] =  9'sd165;
	icos_lut[1238] =  9'sd69;
	qsin_lut[1239] =  9'sd176;
	icos_lut[1239] =  9'sd35;
	qsin_lut[1240] =  9'sd179;
	icos_lut[1240] =  9'sd0;
	qsin_lut[1241] =  9'sd176;
	icos_lut[1241] = -9'sd35;
	qsin_lut[1242] =  9'sd165;
	icos_lut[1242] = -9'sd69;
	qsin_lut[1243] =  9'sd149;
	icos_lut[1243] = -9'sd99;
	qsin_lut[1244] =  9'sd127;
	icos_lut[1244] = -9'sd127;
	qsin_lut[1245] =  9'sd99;
	icos_lut[1245] = -9'sd149;
	qsin_lut[1246] =  9'sd69;
	icos_lut[1246] = -9'sd165;
	qsin_lut[1247] =  9'sd35;
	icos_lut[1247] = -9'sd176;
	qsin_lut[1248] =  9'sd0;
	icos_lut[1248] = -9'sd177;
	qsin_lut[1249] = -9'sd35;
	icos_lut[1249] = -9'sd174;
	qsin_lut[1250] = -9'sd68;
	icos_lut[1250] = -9'sd164;
	qsin_lut[1251] = -9'sd98;
	icos_lut[1251] = -9'sd147;
	qsin_lut[1252] = -9'sd125;
	icos_lut[1252] = -9'sd125;
	qsin_lut[1253] = -9'sd147;
	icos_lut[1253] = -9'sd98;
	qsin_lut[1254] = -9'sd164;
	icos_lut[1254] = -9'sd68;
	qsin_lut[1255] = -9'sd174;
	icos_lut[1255] = -9'sd35;
	qsin_lut[1256] = -9'sd177;
	icos_lut[1256] = -9'sd0;
	qsin_lut[1257] = -9'sd174;
	icos_lut[1257] =  9'sd35;
	qsin_lut[1258] = -9'sd164;
	icos_lut[1258] =  9'sd68;
	qsin_lut[1259] = -9'sd147;
	icos_lut[1259] =  9'sd98;
	qsin_lut[1260] = -9'sd125;
	icos_lut[1260] =  9'sd125;
	qsin_lut[1261] = -9'sd98;
	icos_lut[1261] =  9'sd147;
	qsin_lut[1262] = -9'sd68;
	icos_lut[1262] =  9'sd164;
	qsin_lut[1263] = -9'sd35;
	icos_lut[1263] =  9'sd174;
	qsin_lut[1264] = -9'sd0;
	icos_lut[1264] =  9'sd177;
	qsin_lut[1265] =  9'sd35;
	icos_lut[1265] =  9'sd174;
	qsin_lut[1266] =  9'sd68;
	icos_lut[1266] =  9'sd164;
	qsin_lut[1267] =  9'sd98;
	icos_lut[1267] =  9'sd147;
	qsin_lut[1268] =  9'sd125;
	icos_lut[1268] =  9'sd125;
	qsin_lut[1269] =  9'sd147;
	icos_lut[1269] =  9'sd98;
	qsin_lut[1270] =  9'sd164;
	icos_lut[1270] =  9'sd68;
	qsin_lut[1271] =  9'sd174;
	icos_lut[1271] =  9'sd35;
	qsin_lut[1272] =  9'sd177;
	icos_lut[1272] =  9'sd0;
	qsin_lut[1273] =  9'sd174;
	icos_lut[1273] = -9'sd35;
	qsin_lut[1274] =  9'sd164;
	icos_lut[1274] = -9'sd68;
	qsin_lut[1275] =  9'sd147;
	icos_lut[1275] = -9'sd98;
	qsin_lut[1276] =  9'sd125;
	icos_lut[1276] = -9'sd125;
	qsin_lut[1277] =  9'sd98;
	icos_lut[1277] = -9'sd147;
	qsin_lut[1278] =  9'sd68;
	icos_lut[1278] = -9'sd164;
	qsin_lut[1279] =  9'sd35;
	icos_lut[1279] = -9'sd174;
	qsin_lut[1280] =  9'sd0;
	icos_lut[1280] = -9'sd175;
	qsin_lut[1281] = -9'sd34;
	icos_lut[1281] = -9'sd172;
	qsin_lut[1282] = -9'sd67;
	icos_lut[1282] = -9'sd162;
	qsin_lut[1283] = -9'sd97;
	icos_lut[1283] = -9'sd146;
	qsin_lut[1284] = -9'sd124;
	icos_lut[1284] = -9'sd124;
	qsin_lut[1285] = -9'sd146;
	icos_lut[1285] = -9'sd97;
	qsin_lut[1286] = -9'sd162;
	icos_lut[1286] = -9'sd67;
	qsin_lut[1287] = -9'sd172;
	icos_lut[1287] = -9'sd34;
	qsin_lut[1288] = -9'sd175;
	icos_lut[1288] = -9'sd0;
	qsin_lut[1289] = -9'sd172;
	icos_lut[1289] =  9'sd34;
	qsin_lut[1290] = -9'sd162;
	icos_lut[1290] =  9'sd67;
	qsin_lut[1291] = -9'sd146;
	icos_lut[1291] =  9'sd97;
	qsin_lut[1292] = -9'sd124;
	icos_lut[1292] =  9'sd124;
	qsin_lut[1293] = -9'sd97;
	icos_lut[1293] =  9'sd146;
	qsin_lut[1294] = -9'sd67;
	icos_lut[1294] =  9'sd162;
	qsin_lut[1295] = -9'sd34;
	icos_lut[1295] =  9'sd172;
	qsin_lut[1296] = -9'sd0;
	icos_lut[1296] =  9'sd175;
	qsin_lut[1297] =  9'sd34;
	icos_lut[1297] =  9'sd172;
	qsin_lut[1298] =  9'sd67;
	icos_lut[1298] =  9'sd162;
	qsin_lut[1299] =  9'sd97;
	icos_lut[1299] =  9'sd146;
	qsin_lut[1300] =  9'sd124;
	icos_lut[1300] =  9'sd124;
	qsin_lut[1301] =  9'sd146;
	icos_lut[1301] =  9'sd97;
	qsin_lut[1302] =  9'sd162;
	icos_lut[1302] =  9'sd67;
	qsin_lut[1303] =  9'sd172;
	icos_lut[1303] =  9'sd34;
	qsin_lut[1304] =  9'sd175;
	icos_lut[1304] =  9'sd0;
	qsin_lut[1305] =  9'sd172;
	icos_lut[1305] = -9'sd34;
	qsin_lut[1306] =  9'sd162;
	icos_lut[1306] = -9'sd67;
	qsin_lut[1307] =  9'sd146;
	icos_lut[1307] = -9'sd97;
	qsin_lut[1308] =  9'sd124;
	icos_lut[1308] = -9'sd124;
	qsin_lut[1309] =  9'sd97;
	icos_lut[1309] = -9'sd146;
	qsin_lut[1310] =  9'sd67;
	icos_lut[1310] = -9'sd162;
	qsin_lut[1311] =  9'sd34;
	icos_lut[1311] = -9'sd172;
	qsin_lut[1312] =  9'sd0;
	icos_lut[1312] = -9'sd173;
	qsin_lut[1313] = -9'sd34;
	icos_lut[1313] = -9'sd170;
	qsin_lut[1314] = -9'sd66;
	icos_lut[1314] = -9'sd160;
	qsin_lut[1315] = -9'sd96;
	icos_lut[1315] = -9'sd144;
	qsin_lut[1316] = -9'sd122;
	icos_lut[1316] = -9'sd122;
	qsin_lut[1317] = -9'sd144;
	icos_lut[1317] = -9'sd96;
	qsin_lut[1318] = -9'sd160;
	icos_lut[1318] = -9'sd66;
	qsin_lut[1319] = -9'sd170;
	icos_lut[1319] = -9'sd34;
	qsin_lut[1320] = -9'sd173;
	icos_lut[1320] = -9'sd0;
	qsin_lut[1321] = -9'sd170;
	icos_lut[1321] =  9'sd34;
	qsin_lut[1322] = -9'sd160;
	icos_lut[1322] =  9'sd66;
	qsin_lut[1323] = -9'sd144;
	icos_lut[1323] =  9'sd96;
	qsin_lut[1324] = -9'sd122;
	icos_lut[1324] =  9'sd122;
	qsin_lut[1325] = -9'sd96;
	icos_lut[1325] =  9'sd144;
	qsin_lut[1326] = -9'sd66;
	icos_lut[1326] =  9'sd160;
	qsin_lut[1327] = -9'sd34;
	icos_lut[1327] =  9'sd170;
	qsin_lut[1328] = -9'sd0;
	icos_lut[1328] =  9'sd173;
	qsin_lut[1329] =  9'sd34;
	icos_lut[1329] =  9'sd170;
	qsin_lut[1330] =  9'sd66;
	icos_lut[1330] =  9'sd160;
	qsin_lut[1331] =  9'sd96;
	icos_lut[1331] =  9'sd144;
	qsin_lut[1332] =  9'sd122;
	icos_lut[1332] =  9'sd122;
	qsin_lut[1333] =  9'sd144;
	icos_lut[1333] =  9'sd96;
	qsin_lut[1334] =  9'sd160;
	icos_lut[1334] =  9'sd66;
	qsin_lut[1335] =  9'sd170;
	icos_lut[1335] =  9'sd34;
	qsin_lut[1336] =  9'sd173;
	icos_lut[1336] =  9'sd0;
	qsin_lut[1337] =  9'sd170;
	icos_lut[1337] = -9'sd34;
	qsin_lut[1338] =  9'sd160;
	icos_lut[1338] = -9'sd66;
	qsin_lut[1339] =  9'sd144;
	icos_lut[1339] = -9'sd96;
	qsin_lut[1340] =  9'sd122;
	icos_lut[1340] = -9'sd122;
	qsin_lut[1341] =  9'sd96;
	icos_lut[1341] = -9'sd144;
	qsin_lut[1342] =  9'sd66;
	icos_lut[1342] = -9'sd160;
	qsin_lut[1343] =  9'sd34;
	icos_lut[1343] = -9'sd170;
	qsin_lut[1344] =  9'sd0;
	icos_lut[1344] = -9'sd171;
	qsin_lut[1345] = -9'sd33;
	icos_lut[1345] = -9'sd168;
	qsin_lut[1346] = -9'sd65;
	icos_lut[1346] = -9'sd158;
	qsin_lut[1347] = -9'sd95;
	icos_lut[1347] = -9'sd142;
	qsin_lut[1348] = -9'sd121;
	icos_lut[1348] = -9'sd121;
	qsin_lut[1349] = -9'sd142;
	icos_lut[1349] = -9'sd95;
	qsin_lut[1350] = -9'sd158;
	icos_lut[1350] = -9'sd65;
	qsin_lut[1351] = -9'sd168;
	icos_lut[1351] = -9'sd33;
	qsin_lut[1352] = -9'sd171;
	icos_lut[1352] = -9'sd0;
	qsin_lut[1353] = -9'sd168;
	icos_lut[1353] =  9'sd33;
	qsin_lut[1354] = -9'sd158;
	icos_lut[1354] =  9'sd65;
	qsin_lut[1355] = -9'sd142;
	icos_lut[1355] =  9'sd95;
	qsin_lut[1356] = -9'sd121;
	icos_lut[1356] =  9'sd121;
	qsin_lut[1357] = -9'sd95;
	icos_lut[1357] =  9'sd142;
	qsin_lut[1358] = -9'sd65;
	icos_lut[1358] =  9'sd158;
	qsin_lut[1359] = -9'sd33;
	icos_lut[1359] =  9'sd168;
	qsin_lut[1360] = -9'sd0;
	icos_lut[1360] =  9'sd171;
	qsin_lut[1361] =  9'sd33;
	icos_lut[1361] =  9'sd168;
	qsin_lut[1362] =  9'sd65;
	icos_lut[1362] =  9'sd158;
	qsin_lut[1363] =  9'sd95;
	icos_lut[1363] =  9'sd142;
	qsin_lut[1364] =  9'sd121;
	icos_lut[1364] =  9'sd121;
	qsin_lut[1365] =  9'sd142;
	icos_lut[1365] =  9'sd95;
	qsin_lut[1366] =  9'sd158;
	icos_lut[1366] =  9'sd65;
	qsin_lut[1367] =  9'sd168;
	icos_lut[1367] =  9'sd33;
	qsin_lut[1368] =  9'sd171;
	icos_lut[1368] =  9'sd0;
	qsin_lut[1369] =  9'sd168;
	icos_lut[1369] = -9'sd33;
	qsin_lut[1370] =  9'sd158;
	icos_lut[1370] = -9'sd65;
	qsin_lut[1371] =  9'sd142;
	icos_lut[1371] = -9'sd95;
	qsin_lut[1372] =  9'sd121;
	icos_lut[1372] = -9'sd121;
	qsin_lut[1373] =  9'sd95;
	icos_lut[1373] = -9'sd142;
	qsin_lut[1374] =  9'sd65;
	icos_lut[1374] = -9'sd158;
	qsin_lut[1375] =  9'sd33;
	icos_lut[1375] = -9'sd168;
	qsin_lut[1376] =  9'sd0;
	icos_lut[1376] = -9'sd169;
	qsin_lut[1377] = -9'sd33;
	icos_lut[1377] = -9'sd166;
	qsin_lut[1378] = -9'sd65;
	icos_lut[1378] = -9'sd156;
	qsin_lut[1379] = -9'sd94;
	icos_lut[1379] = -9'sd141;
	qsin_lut[1380] = -9'sd120;
	icos_lut[1380] = -9'sd120;
	qsin_lut[1381] = -9'sd141;
	icos_lut[1381] = -9'sd94;
	qsin_lut[1382] = -9'sd156;
	icos_lut[1382] = -9'sd65;
	qsin_lut[1383] = -9'sd166;
	icos_lut[1383] = -9'sd33;
	qsin_lut[1384] = -9'sd169;
	icos_lut[1384] = -9'sd0;
	qsin_lut[1385] = -9'sd166;
	icos_lut[1385] =  9'sd33;
	qsin_lut[1386] = -9'sd156;
	icos_lut[1386] =  9'sd65;
	qsin_lut[1387] = -9'sd141;
	icos_lut[1387] =  9'sd94;
	qsin_lut[1388] = -9'sd120;
	icos_lut[1388] =  9'sd120;
	qsin_lut[1389] = -9'sd94;
	icos_lut[1389] =  9'sd141;
	qsin_lut[1390] = -9'sd65;
	icos_lut[1390] =  9'sd156;
	qsin_lut[1391] = -9'sd33;
	icos_lut[1391] =  9'sd166;
	qsin_lut[1392] = -9'sd0;
	icos_lut[1392] =  9'sd169;
	qsin_lut[1393] =  9'sd33;
	icos_lut[1393] =  9'sd166;
	qsin_lut[1394] =  9'sd65;
	icos_lut[1394] =  9'sd156;
	qsin_lut[1395] =  9'sd94;
	icos_lut[1395] =  9'sd141;
	qsin_lut[1396] =  9'sd120;
	icos_lut[1396] =  9'sd120;
	qsin_lut[1397] =  9'sd141;
	icos_lut[1397] =  9'sd94;
	qsin_lut[1398] =  9'sd156;
	icos_lut[1398] =  9'sd65;
	qsin_lut[1399] =  9'sd166;
	icos_lut[1399] =  9'sd33;
	qsin_lut[1400] =  9'sd169;
	icos_lut[1400] =  9'sd0;
	qsin_lut[1401] =  9'sd166;
	icos_lut[1401] = -9'sd33;
	qsin_lut[1402] =  9'sd156;
	icos_lut[1402] = -9'sd65;
	qsin_lut[1403] =  9'sd141;
	icos_lut[1403] = -9'sd94;
	qsin_lut[1404] =  9'sd120;
	icos_lut[1404] = -9'sd120;
	qsin_lut[1405] =  9'sd94;
	icos_lut[1405] = -9'sd141;
	qsin_lut[1406] =  9'sd65;
	icos_lut[1406] = -9'sd156;
	qsin_lut[1407] =  9'sd33;
	icos_lut[1407] = -9'sd166;
	qsin_lut[1408] =  9'sd0;
	icos_lut[1408] = -9'sd167;
	qsin_lut[1409] = -9'sd33;
	icos_lut[1409] = -9'sd164;
	qsin_lut[1410] = -9'sd64;
	icos_lut[1410] = -9'sd154;
	qsin_lut[1411] = -9'sd93;
	icos_lut[1411] = -9'sd139;
	qsin_lut[1412] = -9'sd118;
	icos_lut[1412] = -9'sd118;
	qsin_lut[1413] = -9'sd139;
	icos_lut[1413] = -9'sd93;
	qsin_lut[1414] = -9'sd154;
	icos_lut[1414] = -9'sd64;
	qsin_lut[1415] = -9'sd164;
	icos_lut[1415] = -9'sd33;
	qsin_lut[1416] = -9'sd167;
	icos_lut[1416] = -9'sd0;
	qsin_lut[1417] = -9'sd164;
	icos_lut[1417] =  9'sd33;
	qsin_lut[1418] = -9'sd154;
	icos_lut[1418] =  9'sd64;
	qsin_lut[1419] = -9'sd139;
	icos_lut[1419] =  9'sd93;
	qsin_lut[1420] = -9'sd118;
	icos_lut[1420] =  9'sd118;
	qsin_lut[1421] = -9'sd93;
	icos_lut[1421] =  9'sd139;
	qsin_lut[1422] = -9'sd64;
	icos_lut[1422] =  9'sd154;
	qsin_lut[1423] = -9'sd33;
	icos_lut[1423] =  9'sd164;
	qsin_lut[1424] = -9'sd0;
	icos_lut[1424] =  9'sd167;
	qsin_lut[1425] =  9'sd33;
	icos_lut[1425] =  9'sd164;
	qsin_lut[1426] =  9'sd64;
	icos_lut[1426] =  9'sd154;
	qsin_lut[1427] =  9'sd93;
	icos_lut[1427] =  9'sd139;
	qsin_lut[1428] =  9'sd118;
	icos_lut[1428] =  9'sd118;
	qsin_lut[1429] =  9'sd139;
	icos_lut[1429] =  9'sd93;
	qsin_lut[1430] =  9'sd154;
	icos_lut[1430] =  9'sd64;
	qsin_lut[1431] =  9'sd164;
	icos_lut[1431] =  9'sd33;
	qsin_lut[1432] =  9'sd167;
	icos_lut[1432] =  9'sd0;
	qsin_lut[1433] =  9'sd164;
	icos_lut[1433] = -9'sd33;
	qsin_lut[1434] =  9'sd154;
	icos_lut[1434] = -9'sd64;
	qsin_lut[1435] =  9'sd139;
	icos_lut[1435] = -9'sd93;
	qsin_lut[1436] =  9'sd118;
	icos_lut[1436] = -9'sd118;
	qsin_lut[1437] =  9'sd93;
	icos_lut[1437] = -9'sd139;
	qsin_lut[1438] =  9'sd64;
	icos_lut[1438] = -9'sd154;
	qsin_lut[1439] =  9'sd33;
	icos_lut[1439] = -9'sd164;
	qsin_lut[1440] =  9'sd0;
	icos_lut[1440] = -9'sd165;
	qsin_lut[1441] = -9'sd32;
	icos_lut[1441] = -9'sd162;
	qsin_lut[1442] = -9'sd63;
	icos_lut[1442] = -9'sd152;
	qsin_lut[1443] = -9'sd92;
	icos_lut[1443] = -9'sd137;
	qsin_lut[1444] = -9'sd117;
	icos_lut[1444] = -9'sd117;
	qsin_lut[1445] = -9'sd137;
	icos_lut[1445] = -9'sd92;
	qsin_lut[1446] = -9'sd152;
	icos_lut[1446] = -9'sd63;
	qsin_lut[1447] = -9'sd162;
	icos_lut[1447] = -9'sd32;
	qsin_lut[1448] = -9'sd165;
	icos_lut[1448] = -9'sd0;
	qsin_lut[1449] = -9'sd162;
	icos_lut[1449] =  9'sd32;
	qsin_lut[1450] = -9'sd152;
	icos_lut[1450] =  9'sd63;
	qsin_lut[1451] = -9'sd137;
	icos_lut[1451] =  9'sd92;
	qsin_lut[1452] = -9'sd117;
	icos_lut[1452] =  9'sd117;
	qsin_lut[1453] = -9'sd92;
	icos_lut[1453] =  9'sd137;
	qsin_lut[1454] = -9'sd63;
	icos_lut[1454] =  9'sd152;
	qsin_lut[1455] = -9'sd32;
	icos_lut[1455] =  9'sd162;
	qsin_lut[1456] = -9'sd0;
	icos_lut[1456] =  9'sd165;
	qsin_lut[1457] =  9'sd32;
	icos_lut[1457] =  9'sd162;
	qsin_lut[1458] =  9'sd63;
	icos_lut[1458] =  9'sd152;
	qsin_lut[1459] =  9'sd92;
	icos_lut[1459] =  9'sd137;
	qsin_lut[1460] =  9'sd117;
	icos_lut[1460] =  9'sd117;
	qsin_lut[1461] =  9'sd137;
	icos_lut[1461] =  9'sd92;
	qsin_lut[1462] =  9'sd152;
	icos_lut[1462] =  9'sd63;
	qsin_lut[1463] =  9'sd162;
	icos_lut[1463] =  9'sd32;
	qsin_lut[1464] =  9'sd165;
	icos_lut[1464] =  9'sd0;
	qsin_lut[1465] =  9'sd162;
	icos_lut[1465] = -9'sd32;
	qsin_lut[1466] =  9'sd152;
	icos_lut[1466] = -9'sd63;
	qsin_lut[1467] =  9'sd137;
	icos_lut[1467] = -9'sd92;
	qsin_lut[1468] =  9'sd117;
	icos_lut[1468] = -9'sd117;
	qsin_lut[1469] =  9'sd92;
	icos_lut[1469] = -9'sd137;
	qsin_lut[1470] =  9'sd63;
	icos_lut[1470] = -9'sd152;
	qsin_lut[1471] =  9'sd32;
	icos_lut[1471] = -9'sd162;
	qsin_lut[1472] =  9'sd0;
	icos_lut[1472] = -9'sd163;
	qsin_lut[1473] = -9'sd32;
	icos_lut[1473] = -9'sd160;
	qsin_lut[1474] = -9'sd62;
	icos_lut[1474] = -9'sd151;
	qsin_lut[1475] = -9'sd91;
	icos_lut[1475] = -9'sd136;
	qsin_lut[1476] = -9'sd115;
	icos_lut[1476] = -9'sd115;
	qsin_lut[1477] = -9'sd136;
	icos_lut[1477] = -9'sd91;
	qsin_lut[1478] = -9'sd151;
	icos_lut[1478] = -9'sd62;
	qsin_lut[1479] = -9'sd160;
	icos_lut[1479] = -9'sd32;
	qsin_lut[1480] = -9'sd163;
	icos_lut[1480] = -9'sd0;
	qsin_lut[1481] = -9'sd160;
	icos_lut[1481] =  9'sd32;
	qsin_lut[1482] = -9'sd151;
	icos_lut[1482] =  9'sd62;
	qsin_lut[1483] = -9'sd136;
	icos_lut[1483] =  9'sd91;
	qsin_lut[1484] = -9'sd115;
	icos_lut[1484] =  9'sd115;
	qsin_lut[1485] = -9'sd91;
	icos_lut[1485] =  9'sd136;
	qsin_lut[1486] = -9'sd62;
	icos_lut[1486] =  9'sd151;
	qsin_lut[1487] = -9'sd32;
	icos_lut[1487] =  9'sd160;
	qsin_lut[1488] = -9'sd0;
	icos_lut[1488] =  9'sd163;
	qsin_lut[1489] =  9'sd32;
	icos_lut[1489] =  9'sd160;
	qsin_lut[1490] =  9'sd62;
	icos_lut[1490] =  9'sd151;
	qsin_lut[1491] =  9'sd91;
	icos_lut[1491] =  9'sd136;
	qsin_lut[1492] =  9'sd115;
	icos_lut[1492] =  9'sd115;
	qsin_lut[1493] =  9'sd136;
	icos_lut[1493] =  9'sd91;
	qsin_lut[1494] =  9'sd151;
	icos_lut[1494] =  9'sd62;
	qsin_lut[1495] =  9'sd160;
	icos_lut[1495] =  9'sd32;
	qsin_lut[1496] =  9'sd163;
	icos_lut[1496] =  9'sd0;
	qsin_lut[1497] =  9'sd160;
	icos_lut[1497] = -9'sd32;
	qsin_lut[1498] =  9'sd151;
	icos_lut[1498] = -9'sd62;
	qsin_lut[1499] =  9'sd136;
	icos_lut[1499] = -9'sd91;
	qsin_lut[1500] =  9'sd115;
	icos_lut[1500] = -9'sd115;
	qsin_lut[1501] =  9'sd91;
	icos_lut[1501] = -9'sd136;
	qsin_lut[1502] =  9'sd62;
	icos_lut[1502] = -9'sd151;
	qsin_lut[1503] =  9'sd32;
	icos_lut[1503] = -9'sd160;
	qsin_lut[1504] =  9'sd0;
	icos_lut[1504] = -9'sd161;
	qsin_lut[1505] = -9'sd31;
	icos_lut[1505] = -9'sd158;
	qsin_lut[1506] = -9'sd62;
	icos_lut[1506] = -9'sd149;
	qsin_lut[1507] = -9'sd89;
	icos_lut[1507] = -9'sd134;
	qsin_lut[1508] = -9'sd114;
	icos_lut[1508] = -9'sd114;
	qsin_lut[1509] = -9'sd134;
	icos_lut[1509] = -9'sd89;
	qsin_lut[1510] = -9'sd149;
	icos_lut[1510] = -9'sd62;
	qsin_lut[1511] = -9'sd158;
	icos_lut[1511] = -9'sd31;
	qsin_lut[1512] = -9'sd161;
	icos_lut[1512] = -9'sd0;
	qsin_lut[1513] = -9'sd158;
	icos_lut[1513] =  9'sd31;
	qsin_lut[1514] = -9'sd149;
	icos_lut[1514] =  9'sd62;
	qsin_lut[1515] = -9'sd134;
	icos_lut[1515] =  9'sd89;
	qsin_lut[1516] = -9'sd114;
	icos_lut[1516] =  9'sd114;
	qsin_lut[1517] = -9'sd89;
	icos_lut[1517] =  9'sd134;
	qsin_lut[1518] = -9'sd62;
	icos_lut[1518] =  9'sd149;
	qsin_lut[1519] = -9'sd31;
	icos_lut[1519] =  9'sd158;
	qsin_lut[1520] = -9'sd0;
	icos_lut[1520] =  9'sd161;
	qsin_lut[1521] =  9'sd31;
	icos_lut[1521] =  9'sd158;
	qsin_lut[1522] =  9'sd62;
	icos_lut[1522] =  9'sd149;
	qsin_lut[1523] =  9'sd89;
	icos_lut[1523] =  9'sd134;
	qsin_lut[1524] =  9'sd114;
	icos_lut[1524] =  9'sd114;
	qsin_lut[1525] =  9'sd134;
	icos_lut[1525] =  9'sd89;
	qsin_lut[1526] =  9'sd149;
	icos_lut[1526] =  9'sd62;
	qsin_lut[1527] =  9'sd158;
	icos_lut[1527] =  9'sd31;
	qsin_lut[1528] =  9'sd161;
	icos_lut[1528] =  9'sd0;
	qsin_lut[1529] =  9'sd158;
	icos_lut[1529] = -9'sd31;
	qsin_lut[1530] =  9'sd149;
	icos_lut[1530] = -9'sd62;
	qsin_lut[1531] =  9'sd134;
	icos_lut[1531] = -9'sd89;
	qsin_lut[1532] =  9'sd114;
	icos_lut[1532] = -9'sd114;
	qsin_lut[1533] =  9'sd89;
	icos_lut[1533] = -9'sd134;
	qsin_lut[1534] =  9'sd62;
	icos_lut[1534] = -9'sd149;
	qsin_lut[1535] =  9'sd31;
	icos_lut[1535] = -9'sd158;
	qsin_lut[1536] =  9'sd0;
	icos_lut[1536] = -9'sd159;
	qsin_lut[1537] = -9'sd31;
	icos_lut[1537] = -9'sd156;
	qsin_lut[1538] = -9'sd61;
	icos_lut[1538] = -9'sd147;
	qsin_lut[1539] = -9'sd88;
	icos_lut[1539] = -9'sd132;
	qsin_lut[1540] = -9'sd112;
	icos_lut[1540] = -9'sd112;
	qsin_lut[1541] = -9'sd132;
	icos_lut[1541] = -9'sd88;
	qsin_lut[1542] = -9'sd147;
	icos_lut[1542] = -9'sd61;
	qsin_lut[1543] = -9'sd156;
	icos_lut[1543] = -9'sd31;
	qsin_lut[1544] = -9'sd159;
	icos_lut[1544] = -9'sd0;
	qsin_lut[1545] = -9'sd156;
	icos_lut[1545] =  9'sd31;
	qsin_lut[1546] = -9'sd147;
	icos_lut[1546] =  9'sd61;
	qsin_lut[1547] = -9'sd132;
	icos_lut[1547] =  9'sd88;
	qsin_lut[1548] = -9'sd112;
	icos_lut[1548] =  9'sd112;
	qsin_lut[1549] = -9'sd88;
	icos_lut[1549] =  9'sd132;
	qsin_lut[1550] = -9'sd61;
	icos_lut[1550] =  9'sd147;
	qsin_lut[1551] = -9'sd31;
	icos_lut[1551] =  9'sd156;
	qsin_lut[1552] = -9'sd0;
	icos_lut[1552] =  9'sd159;
	qsin_lut[1553] =  9'sd31;
	icos_lut[1553] =  9'sd156;
	qsin_lut[1554] =  9'sd61;
	icos_lut[1554] =  9'sd147;
	qsin_lut[1555] =  9'sd88;
	icos_lut[1555] =  9'sd132;
	qsin_lut[1556] =  9'sd112;
	icos_lut[1556] =  9'sd112;
	qsin_lut[1557] =  9'sd132;
	icos_lut[1557] =  9'sd88;
	qsin_lut[1558] =  9'sd147;
	icos_lut[1558] =  9'sd61;
	qsin_lut[1559] =  9'sd156;
	icos_lut[1559] =  9'sd31;
	qsin_lut[1560] =  9'sd159;
	icos_lut[1560] =  9'sd0;
	qsin_lut[1561] =  9'sd156;
	icos_lut[1561] = -9'sd31;
	qsin_lut[1562] =  9'sd147;
	icos_lut[1562] = -9'sd61;
	qsin_lut[1563] =  9'sd132;
	icos_lut[1563] = -9'sd88;
	qsin_lut[1564] =  9'sd112;
	icos_lut[1564] = -9'sd112;
	qsin_lut[1565] =  9'sd88;
	icos_lut[1565] = -9'sd132;
	qsin_lut[1566] =  9'sd61;
	icos_lut[1566] = -9'sd147;
	qsin_lut[1567] =  9'sd31;
	icos_lut[1567] = -9'sd156;
	qsin_lut[1568] =  9'sd0;
	icos_lut[1568] = -9'sd157;
	qsin_lut[1569] = -9'sd31;
	icos_lut[1569] = -9'sd154;
	qsin_lut[1570] = -9'sd60;
	icos_lut[1570] = -9'sd145;
	qsin_lut[1571] = -9'sd87;
	icos_lut[1571] = -9'sd131;
	qsin_lut[1572] = -9'sd111;
	icos_lut[1572] = -9'sd111;
	qsin_lut[1573] = -9'sd131;
	icos_lut[1573] = -9'sd87;
	qsin_lut[1574] = -9'sd145;
	icos_lut[1574] = -9'sd60;
	qsin_lut[1575] = -9'sd154;
	icos_lut[1575] = -9'sd31;
	qsin_lut[1576] = -9'sd157;
	icos_lut[1576] = -9'sd0;
	qsin_lut[1577] = -9'sd154;
	icos_lut[1577] =  9'sd31;
	qsin_lut[1578] = -9'sd145;
	icos_lut[1578] =  9'sd60;
	qsin_lut[1579] = -9'sd131;
	icos_lut[1579] =  9'sd87;
	qsin_lut[1580] = -9'sd111;
	icos_lut[1580] =  9'sd111;
	qsin_lut[1581] = -9'sd87;
	icos_lut[1581] =  9'sd131;
	qsin_lut[1582] = -9'sd60;
	icos_lut[1582] =  9'sd145;
	qsin_lut[1583] = -9'sd31;
	icos_lut[1583] =  9'sd154;
	qsin_lut[1584] = -9'sd0;
	icos_lut[1584] =  9'sd157;
	qsin_lut[1585] =  9'sd31;
	icos_lut[1585] =  9'sd154;
	qsin_lut[1586] =  9'sd60;
	icos_lut[1586] =  9'sd145;
	qsin_lut[1587] =  9'sd87;
	icos_lut[1587] =  9'sd131;
	qsin_lut[1588] =  9'sd111;
	icos_lut[1588] =  9'sd111;
	qsin_lut[1589] =  9'sd131;
	icos_lut[1589] =  9'sd87;
	qsin_lut[1590] =  9'sd145;
	icos_lut[1590] =  9'sd60;
	qsin_lut[1591] =  9'sd154;
	icos_lut[1591] =  9'sd31;
	qsin_lut[1592] =  9'sd157;
	icos_lut[1592] =  9'sd0;
	qsin_lut[1593] =  9'sd154;
	icos_lut[1593] = -9'sd31;
	qsin_lut[1594] =  9'sd145;
	icos_lut[1594] = -9'sd60;
	qsin_lut[1595] =  9'sd131;
	icos_lut[1595] = -9'sd87;
	qsin_lut[1596] =  9'sd111;
	icos_lut[1596] = -9'sd111;
	qsin_lut[1597] =  9'sd87;
	icos_lut[1597] = -9'sd131;
	qsin_lut[1598] =  9'sd60;
	icos_lut[1598] = -9'sd145;
	qsin_lut[1599] =  9'sd31;
	icos_lut[1599] = -9'sd154;
	qsin_lut[1600] =  9'sd0;
	icos_lut[1600] = -9'sd155;
	qsin_lut[1601] = -9'sd30;
	icos_lut[1601] = -9'sd152;
	qsin_lut[1602] = -9'sd59;
	icos_lut[1602] = -9'sd143;
	qsin_lut[1603] = -9'sd86;
	icos_lut[1603] = -9'sd129;
	qsin_lut[1604] = -9'sd110;
	icos_lut[1604] = -9'sd110;
	qsin_lut[1605] = -9'sd129;
	icos_lut[1605] = -9'sd86;
	qsin_lut[1606] = -9'sd143;
	icos_lut[1606] = -9'sd59;
	qsin_lut[1607] = -9'sd152;
	icos_lut[1607] = -9'sd30;
	qsin_lut[1608] = -9'sd155;
	icos_lut[1608] = -9'sd0;
	qsin_lut[1609] = -9'sd152;
	icos_lut[1609] =  9'sd30;
	qsin_lut[1610] = -9'sd143;
	icos_lut[1610] =  9'sd59;
	qsin_lut[1611] = -9'sd129;
	icos_lut[1611] =  9'sd86;
	qsin_lut[1612] = -9'sd110;
	icos_lut[1612] =  9'sd110;
	qsin_lut[1613] = -9'sd86;
	icos_lut[1613] =  9'sd129;
	qsin_lut[1614] = -9'sd59;
	icos_lut[1614] =  9'sd143;
	qsin_lut[1615] = -9'sd30;
	icos_lut[1615] =  9'sd152;
	qsin_lut[1616] = -9'sd0;
	icos_lut[1616] =  9'sd155;
	qsin_lut[1617] =  9'sd30;
	icos_lut[1617] =  9'sd152;
	qsin_lut[1618] =  9'sd59;
	icos_lut[1618] =  9'sd143;
	qsin_lut[1619] =  9'sd86;
	icos_lut[1619] =  9'sd129;
	qsin_lut[1620] =  9'sd110;
	icos_lut[1620] =  9'sd110;
	qsin_lut[1621] =  9'sd129;
	icos_lut[1621] =  9'sd86;
	qsin_lut[1622] =  9'sd143;
	icos_lut[1622] =  9'sd59;
	qsin_lut[1623] =  9'sd152;
	icos_lut[1623] =  9'sd30;
	qsin_lut[1624] =  9'sd155;
	icos_lut[1624] =  9'sd0;
	qsin_lut[1625] =  9'sd152;
	icos_lut[1625] = -9'sd30;
	qsin_lut[1626] =  9'sd143;
	icos_lut[1626] = -9'sd59;
	qsin_lut[1627] =  9'sd129;
	icos_lut[1627] = -9'sd86;
	qsin_lut[1628] =  9'sd110;
	icos_lut[1628] = -9'sd110;
	qsin_lut[1629] =  9'sd86;
	icos_lut[1629] = -9'sd129;
	qsin_lut[1630] =  9'sd59;
	icos_lut[1630] = -9'sd143;
	qsin_lut[1631] =  9'sd30;
	icos_lut[1631] = -9'sd152;
	qsin_lut[1632] =  9'sd0;
	icos_lut[1632] = -9'sd153;
	qsin_lut[1633] = -9'sd30;
	icos_lut[1633] = -9'sd150;
	qsin_lut[1634] = -9'sd59;
	icos_lut[1634] = -9'sd141;
	qsin_lut[1635] = -9'sd85;
	icos_lut[1635] = -9'sd127;
	qsin_lut[1636] = -9'sd108;
	icos_lut[1636] = -9'sd108;
	qsin_lut[1637] = -9'sd127;
	icos_lut[1637] = -9'sd85;
	qsin_lut[1638] = -9'sd141;
	icos_lut[1638] = -9'sd59;
	qsin_lut[1639] = -9'sd150;
	icos_lut[1639] = -9'sd30;
	qsin_lut[1640] = -9'sd153;
	icos_lut[1640] = -9'sd0;
	qsin_lut[1641] = -9'sd150;
	icos_lut[1641] =  9'sd30;
	qsin_lut[1642] = -9'sd141;
	icos_lut[1642] =  9'sd59;
	qsin_lut[1643] = -9'sd127;
	icos_lut[1643] =  9'sd85;
	qsin_lut[1644] = -9'sd108;
	icos_lut[1644] =  9'sd108;
	qsin_lut[1645] = -9'sd85;
	icos_lut[1645] =  9'sd127;
	qsin_lut[1646] = -9'sd59;
	icos_lut[1646] =  9'sd141;
	qsin_lut[1647] = -9'sd30;
	icos_lut[1647] =  9'sd150;
	qsin_lut[1648] = -9'sd0;
	icos_lut[1648] =  9'sd153;
	qsin_lut[1649] =  9'sd30;
	icos_lut[1649] =  9'sd150;
	qsin_lut[1650] =  9'sd59;
	icos_lut[1650] =  9'sd141;
	qsin_lut[1651] =  9'sd85;
	icos_lut[1651] =  9'sd127;
	qsin_lut[1652] =  9'sd108;
	icos_lut[1652] =  9'sd108;
	qsin_lut[1653] =  9'sd127;
	icos_lut[1653] =  9'sd85;
	qsin_lut[1654] =  9'sd141;
	icos_lut[1654] =  9'sd59;
	qsin_lut[1655] =  9'sd150;
	icos_lut[1655] =  9'sd30;
	qsin_lut[1656] =  9'sd153;
	icos_lut[1656] =  9'sd0;
	qsin_lut[1657] =  9'sd150;
	icos_lut[1657] = -9'sd30;
	qsin_lut[1658] =  9'sd141;
	icos_lut[1658] = -9'sd59;
	qsin_lut[1659] =  9'sd127;
	icos_lut[1659] = -9'sd85;
	qsin_lut[1660] =  9'sd108;
	icos_lut[1660] = -9'sd108;
	qsin_lut[1661] =  9'sd85;
	icos_lut[1661] = -9'sd127;
	qsin_lut[1662] =  9'sd59;
	icos_lut[1662] = -9'sd141;
	qsin_lut[1663] =  9'sd30;
	icos_lut[1663] = -9'sd150;
	qsin_lut[1664] =  9'sd0;
	icos_lut[1664] = -9'sd151;
	qsin_lut[1665] = -9'sd29;
	icos_lut[1665] = -9'sd148;
	qsin_lut[1666] = -9'sd58;
	icos_lut[1666] = -9'sd140;
	qsin_lut[1667] = -9'sd84;
	icos_lut[1667] = -9'sd126;
	qsin_lut[1668] = -9'sd107;
	icos_lut[1668] = -9'sd107;
	qsin_lut[1669] = -9'sd126;
	icos_lut[1669] = -9'sd84;
	qsin_lut[1670] = -9'sd140;
	icos_lut[1670] = -9'sd58;
	qsin_lut[1671] = -9'sd148;
	icos_lut[1671] = -9'sd29;
	qsin_lut[1672] = -9'sd151;
	icos_lut[1672] = -9'sd0;
	qsin_lut[1673] = -9'sd148;
	icos_lut[1673] =  9'sd29;
	qsin_lut[1674] = -9'sd140;
	icos_lut[1674] =  9'sd58;
	qsin_lut[1675] = -9'sd126;
	icos_lut[1675] =  9'sd84;
	qsin_lut[1676] = -9'sd107;
	icos_lut[1676] =  9'sd107;
	qsin_lut[1677] = -9'sd84;
	icos_lut[1677] =  9'sd126;
	qsin_lut[1678] = -9'sd58;
	icos_lut[1678] =  9'sd140;
	qsin_lut[1679] = -9'sd29;
	icos_lut[1679] =  9'sd148;
	qsin_lut[1680] = -9'sd0;
	icos_lut[1680] =  9'sd151;
	qsin_lut[1681] =  9'sd29;
	icos_lut[1681] =  9'sd148;
	qsin_lut[1682] =  9'sd58;
	icos_lut[1682] =  9'sd140;
	qsin_lut[1683] =  9'sd84;
	icos_lut[1683] =  9'sd126;
	qsin_lut[1684] =  9'sd107;
	icos_lut[1684] =  9'sd107;
	qsin_lut[1685] =  9'sd126;
	icos_lut[1685] =  9'sd84;
	qsin_lut[1686] =  9'sd140;
	icos_lut[1686] =  9'sd58;
	qsin_lut[1687] =  9'sd148;
	icos_lut[1687] =  9'sd29;
	qsin_lut[1688] =  9'sd151;
	icos_lut[1688] =  9'sd0;
	qsin_lut[1689] =  9'sd148;
	icos_lut[1689] = -9'sd29;
	qsin_lut[1690] =  9'sd140;
	icos_lut[1690] = -9'sd58;
	qsin_lut[1691] =  9'sd126;
	icos_lut[1691] = -9'sd84;
	qsin_lut[1692] =  9'sd107;
	icos_lut[1692] = -9'sd107;
	qsin_lut[1693] =  9'sd84;
	icos_lut[1693] = -9'sd126;
	qsin_lut[1694] =  9'sd58;
	icos_lut[1694] = -9'sd140;
	qsin_lut[1695] =  9'sd29;
	icos_lut[1695] = -9'sd148;
	qsin_lut[1696] =  9'sd0;
	icos_lut[1696] = -9'sd149;
	qsin_lut[1697] = -9'sd29;
	icos_lut[1697] = -9'sd146;
	qsin_lut[1698] = -9'sd57;
	icos_lut[1698] = -9'sd138;
	qsin_lut[1699] = -9'sd83;
	icos_lut[1699] = -9'sd124;
	qsin_lut[1700] = -9'sd105;
	icos_lut[1700] = -9'sd105;
	qsin_lut[1701] = -9'sd124;
	icos_lut[1701] = -9'sd83;
	qsin_lut[1702] = -9'sd138;
	icos_lut[1702] = -9'sd57;
	qsin_lut[1703] = -9'sd146;
	icos_lut[1703] = -9'sd29;
	qsin_lut[1704] = -9'sd149;
	icos_lut[1704] = -9'sd0;
	qsin_lut[1705] = -9'sd146;
	icos_lut[1705] =  9'sd29;
	qsin_lut[1706] = -9'sd138;
	icos_lut[1706] =  9'sd57;
	qsin_lut[1707] = -9'sd124;
	icos_lut[1707] =  9'sd83;
	qsin_lut[1708] = -9'sd105;
	icos_lut[1708] =  9'sd105;
	qsin_lut[1709] = -9'sd83;
	icos_lut[1709] =  9'sd124;
	qsin_lut[1710] = -9'sd57;
	icos_lut[1710] =  9'sd138;
	qsin_lut[1711] = -9'sd29;
	icos_lut[1711] =  9'sd146;
	qsin_lut[1712] = -9'sd0;
	icos_lut[1712] =  9'sd149;
	qsin_lut[1713] =  9'sd29;
	icos_lut[1713] =  9'sd146;
	qsin_lut[1714] =  9'sd57;
	icos_lut[1714] =  9'sd138;
	qsin_lut[1715] =  9'sd83;
	icos_lut[1715] =  9'sd124;
	qsin_lut[1716] =  9'sd105;
	icos_lut[1716] =  9'sd105;
	qsin_lut[1717] =  9'sd124;
	icos_lut[1717] =  9'sd83;
	qsin_lut[1718] =  9'sd138;
	icos_lut[1718] =  9'sd57;
	qsin_lut[1719] =  9'sd146;
	icos_lut[1719] =  9'sd29;
	qsin_lut[1720] =  9'sd149;
	icos_lut[1720] =  9'sd0;
	qsin_lut[1721] =  9'sd146;
	icos_lut[1721] = -9'sd29;
	qsin_lut[1722] =  9'sd138;
	icos_lut[1722] = -9'sd57;
	qsin_lut[1723] =  9'sd124;
	icos_lut[1723] = -9'sd83;
	qsin_lut[1724] =  9'sd105;
	icos_lut[1724] = -9'sd105;
	qsin_lut[1725] =  9'sd83;
	icos_lut[1725] = -9'sd124;
	qsin_lut[1726] =  9'sd57;
	icos_lut[1726] = -9'sd138;
	qsin_lut[1727] =  9'sd29;
	icos_lut[1727] = -9'sd146;
	qsin_lut[1728] =  9'sd0;
	icos_lut[1728] = -9'sd147;
	qsin_lut[1729] = -9'sd29;
	icos_lut[1729] = -9'sd144;
	qsin_lut[1730] = -9'sd56;
	icos_lut[1730] = -9'sd136;
	qsin_lut[1731] = -9'sd82;
	icos_lut[1731] = -9'sd122;
	qsin_lut[1732] = -9'sd104;
	icos_lut[1732] = -9'sd104;
	qsin_lut[1733] = -9'sd122;
	icos_lut[1733] = -9'sd82;
	qsin_lut[1734] = -9'sd136;
	icos_lut[1734] = -9'sd56;
	qsin_lut[1735] = -9'sd144;
	icos_lut[1735] = -9'sd29;
	qsin_lut[1736] = -9'sd147;
	icos_lut[1736] = -9'sd0;
	qsin_lut[1737] = -9'sd144;
	icos_lut[1737] =  9'sd29;
	qsin_lut[1738] = -9'sd136;
	icos_lut[1738] =  9'sd56;
	qsin_lut[1739] = -9'sd122;
	icos_lut[1739] =  9'sd82;
	qsin_lut[1740] = -9'sd104;
	icos_lut[1740] =  9'sd104;
	qsin_lut[1741] = -9'sd82;
	icos_lut[1741] =  9'sd122;
	qsin_lut[1742] = -9'sd56;
	icos_lut[1742] =  9'sd136;
	qsin_lut[1743] = -9'sd29;
	icos_lut[1743] =  9'sd144;
	qsin_lut[1744] = -9'sd0;
	icos_lut[1744] =  9'sd147;
	qsin_lut[1745] =  9'sd29;
	icos_lut[1745] =  9'sd144;
	qsin_lut[1746] =  9'sd56;
	icos_lut[1746] =  9'sd136;
	qsin_lut[1747] =  9'sd82;
	icos_lut[1747] =  9'sd122;
	qsin_lut[1748] =  9'sd104;
	icos_lut[1748] =  9'sd104;
	qsin_lut[1749] =  9'sd122;
	icos_lut[1749] =  9'sd82;
	qsin_lut[1750] =  9'sd136;
	icos_lut[1750] =  9'sd56;
	qsin_lut[1751] =  9'sd144;
	icos_lut[1751] =  9'sd29;
	qsin_lut[1752] =  9'sd147;
	icos_lut[1752] =  9'sd0;
	qsin_lut[1753] =  9'sd144;
	icos_lut[1753] = -9'sd29;
	qsin_lut[1754] =  9'sd136;
	icos_lut[1754] = -9'sd56;
	qsin_lut[1755] =  9'sd122;
	icos_lut[1755] = -9'sd82;
	qsin_lut[1756] =  9'sd104;
	icos_lut[1756] = -9'sd104;
	qsin_lut[1757] =  9'sd82;
	icos_lut[1757] = -9'sd122;
	qsin_lut[1758] =  9'sd56;
	icos_lut[1758] = -9'sd136;
	qsin_lut[1759] =  9'sd29;
	icos_lut[1759] = -9'sd144;
	qsin_lut[1760] =  9'sd0;
	icos_lut[1760] = -9'sd145;
	qsin_lut[1761] = -9'sd28;
	icos_lut[1761] = -9'sd142;
	qsin_lut[1762] = -9'sd55;
	icos_lut[1762] = -9'sd134;
	qsin_lut[1763] = -9'sd81;
	icos_lut[1763] = -9'sd121;
	qsin_lut[1764] = -9'sd103;
	icos_lut[1764] = -9'sd103;
	qsin_lut[1765] = -9'sd121;
	icos_lut[1765] = -9'sd81;
	qsin_lut[1766] = -9'sd134;
	icos_lut[1766] = -9'sd55;
	qsin_lut[1767] = -9'sd142;
	icos_lut[1767] = -9'sd28;
	qsin_lut[1768] = -9'sd145;
	icos_lut[1768] = -9'sd0;
	qsin_lut[1769] = -9'sd142;
	icos_lut[1769] =  9'sd28;
	qsin_lut[1770] = -9'sd134;
	icos_lut[1770] =  9'sd55;
	qsin_lut[1771] = -9'sd121;
	icos_lut[1771] =  9'sd81;
	qsin_lut[1772] = -9'sd103;
	icos_lut[1772] =  9'sd103;
	qsin_lut[1773] = -9'sd81;
	icos_lut[1773] =  9'sd121;
	qsin_lut[1774] = -9'sd55;
	icos_lut[1774] =  9'sd134;
	qsin_lut[1775] = -9'sd28;
	icos_lut[1775] =  9'sd142;
	qsin_lut[1776] = -9'sd0;
	icos_lut[1776] =  9'sd145;
	qsin_lut[1777] =  9'sd28;
	icos_lut[1777] =  9'sd142;
	qsin_lut[1778] =  9'sd55;
	icos_lut[1778] =  9'sd134;
	qsin_lut[1779] =  9'sd81;
	icos_lut[1779] =  9'sd121;
	qsin_lut[1780] =  9'sd103;
	icos_lut[1780] =  9'sd103;
	qsin_lut[1781] =  9'sd121;
	icos_lut[1781] =  9'sd81;
	qsin_lut[1782] =  9'sd134;
	icos_lut[1782] =  9'sd55;
	qsin_lut[1783] =  9'sd142;
	icos_lut[1783] =  9'sd28;
	qsin_lut[1784] =  9'sd145;
	icos_lut[1784] =  9'sd0;
	qsin_lut[1785] =  9'sd142;
	icos_lut[1785] = -9'sd28;
	qsin_lut[1786] =  9'sd134;
	icos_lut[1786] = -9'sd55;
	qsin_lut[1787] =  9'sd121;
	icos_lut[1787] = -9'sd81;
	qsin_lut[1788] =  9'sd103;
	icos_lut[1788] = -9'sd103;
	qsin_lut[1789] =  9'sd81;
	icos_lut[1789] = -9'sd121;
	qsin_lut[1790] =  9'sd55;
	icos_lut[1790] = -9'sd134;
	qsin_lut[1791] =  9'sd28;
	icos_lut[1791] = -9'sd142;
	qsin_lut[1792] =  9'sd0;
	icos_lut[1792] = -9'sd143;
	qsin_lut[1793] = -9'sd28;
	icos_lut[1793] = -9'sd140;
	qsin_lut[1794] = -9'sd55;
	icos_lut[1794] = -9'sd132;
	qsin_lut[1795] = -9'sd79;
	icos_lut[1795] = -9'sd119;
	qsin_lut[1796] = -9'sd101;
	icos_lut[1796] = -9'sd101;
	qsin_lut[1797] = -9'sd119;
	icos_lut[1797] = -9'sd79;
	qsin_lut[1798] = -9'sd132;
	icos_lut[1798] = -9'sd55;
	qsin_lut[1799] = -9'sd140;
	icos_lut[1799] = -9'sd28;
	qsin_lut[1800] = -9'sd143;
	icos_lut[1800] = -9'sd0;
	qsin_lut[1801] = -9'sd140;
	icos_lut[1801] =  9'sd28;
	qsin_lut[1802] = -9'sd132;
	icos_lut[1802] =  9'sd55;
	qsin_lut[1803] = -9'sd119;
	icos_lut[1803] =  9'sd79;
	qsin_lut[1804] = -9'sd101;
	icos_lut[1804] =  9'sd101;
	qsin_lut[1805] = -9'sd79;
	icos_lut[1805] =  9'sd119;
	qsin_lut[1806] = -9'sd55;
	icos_lut[1806] =  9'sd132;
	qsin_lut[1807] = -9'sd28;
	icos_lut[1807] =  9'sd140;
	qsin_lut[1808] = -9'sd0;
	icos_lut[1808] =  9'sd143;
	qsin_lut[1809] =  9'sd28;
	icos_lut[1809] =  9'sd140;
	qsin_lut[1810] =  9'sd55;
	icos_lut[1810] =  9'sd132;
	qsin_lut[1811] =  9'sd79;
	icos_lut[1811] =  9'sd119;
	qsin_lut[1812] =  9'sd101;
	icos_lut[1812] =  9'sd101;
	qsin_lut[1813] =  9'sd119;
	icos_lut[1813] =  9'sd79;
	qsin_lut[1814] =  9'sd132;
	icos_lut[1814] =  9'sd55;
	qsin_lut[1815] =  9'sd140;
	icos_lut[1815] =  9'sd28;
	qsin_lut[1816] =  9'sd143;
	icos_lut[1816] =  9'sd0;
	qsin_lut[1817] =  9'sd140;
	icos_lut[1817] = -9'sd28;
	qsin_lut[1818] =  9'sd132;
	icos_lut[1818] = -9'sd55;
	qsin_lut[1819] =  9'sd119;
	icos_lut[1819] = -9'sd79;
	qsin_lut[1820] =  9'sd101;
	icos_lut[1820] = -9'sd101;
	qsin_lut[1821] =  9'sd79;
	icos_lut[1821] = -9'sd119;
	qsin_lut[1822] =  9'sd55;
	icos_lut[1822] = -9'sd132;
	qsin_lut[1823] =  9'sd28;
	icos_lut[1823] = -9'sd140;
	qsin_lut[1824] =  9'sd0;
	icos_lut[1824] = -9'sd141;
	qsin_lut[1825] = -9'sd28;
	icos_lut[1825] = -9'sd138;
	qsin_lut[1826] = -9'sd54;
	icos_lut[1826] = -9'sd130;
	qsin_lut[1827] = -9'sd78;
	icos_lut[1827] = -9'sd117;
	qsin_lut[1828] = -9'sd100;
	icos_lut[1828] = -9'sd100;
	qsin_lut[1829] = -9'sd117;
	icos_lut[1829] = -9'sd78;
	qsin_lut[1830] = -9'sd130;
	icos_lut[1830] = -9'sd54;
	qsin_lut[1831] = -9'sd138;
	icos_lut[1831] = -9'sd28;
	qsin_lut[1832] = -9'sd141;
	icos_lut[1832] = -9'sd0;
	qsin_lut[1833] = -9'sd138;
	icos_lut[1833] =  9'sd28;
	qsin_lut[1834] = -9'sd130;
	icos_lut[1834] =  9'sd54;
	qsin_lut[1835] = -9'sd117;
	icos_lut[1835] =  9'sd78;
	qsin_lut[1836] = -9'sd100;
	icos_lut[1836] =  9'sd100;
	qsin_lut[1837] = -9'sd78;
	icos_lut[1837] =  9'sd117;
	qsin_lut[1838] = -9'sd54;
	icos_lut[1838] =  9'sd130;
	qsin_lut[1839] = -9'sd28;
	icos_lut[1839] =  9'sd138;
	qsin_lut[1840] = -9'sd0;
	icos_lut[1840] =  9'sd141;
	qsin_lut[1841] =  9'sd28;
	icos_lut[1841] =  9'sd138;
	qsin_lut[1842] =  9'sd54;
	icos_lut[1842] =  9'sd130;
	qsin_lut[1843] =  9'sd78;
	icos_lut[1843] =  9'sd117;
	qsin_lut[1844] =  9'sd100;
	icos_lut[1844] =  9'sd100;
	qsin_lut[1845] =  9'sd117;
	icos_lut[1845] =  9'sd78;
	qsin_lut[1846] =  9'sd130;
	icos_lut[1846] =  9'sd54;
	qsin_lut[1847] =  9'sd138;
	icos_lut[1847] =  9'sd28;
	qsin_lut[1848] =  9'sd141;
	icos_lut[1848] =  9'sd0;
	qsin_lut[1849] =  9'sd138;
	icos_lut[1849] = -9'sd28;
	qsin_lut[1850] =  9'sd130;
	icos_lut[1850] = -9'sd54;
	qsin_lut[1851] =  9'sd117;
	icos_lut[1851] = -9'sd78;
	qsin_lut[1852] =  9'sd100;
	icos_lut[1852] = -9'sd100;
	qsin_lut[1853] =  9'sd78;
	icos_lut[1853] = -9'sd117;
	qsin_lut[1854] =  9'sd54;
	icos_lut[1854] = -9'sd130;
	qsin_lut[1855] =  9'sd28;
	icos_lut[1855] = -9'sd138;
	qsin_lut[1856] =  9'sd0;
	icos_lut[1856] = -9'sd139;
	qsin_lut[1857] = -9'sd27;
	icos_lut[1857] = -9'sd136;
	qsin_lut[1858] = -9'sd53;
	icos_lut[1858] = -9'sd128;
	qsin_lut[1859] = -9'sd77;
	icos_lut[1859] = -9'sd116;
	qsin_lut[1860] = -9'sd98;
	icos_lut[1860] = -9'sd98;
	qsin_lut[1861] = -9'sd116;
	icos_lut[1861] = -9'sd77;
	qsin_lut[1862] = -9'sd128;
	icos_lut[1862] = -9'sd53;
	qsin_lut[1863] = -9'sd136;
	icos_lut[1863] = -9'sd27;
	qsin_lut[1864] = -9'sd139;
	icos_lut[1864] = -9'sd0;
	qsin_lut[1865] = -9'sd136;
	icos_lut[1865] =  9'sd27;
	qsin_lut[1866] = -9'sd128;
	icos_lut[1866] =  9'sd53;
	qsin_lut[1867] = -9'sd116;
	icos_lut[1867] =  9'sd77;
	qsin_lut[1868] = -9'sd98;
	icos_lut[1868] =  9'sd98;
	qsin_lut[1869] = -9'sd77;
	icos_lut[1869] =  9'sd116;
	qsin_lut[1870] = -9'sd53;
	icos_lut[1870] =  9'sd128;
	qsin_lut[1871] = -9'sd27;
	icos_lut[1871] =  9'sd136;
	qsin_lut[1872] = -9'sd0;
	icos_lut[1872] =  9'sd139;
	qsin_lut[1873] =  9'sd27;
	icos_lut[1873] =  9'sd136;
	qsin_lut[1874] =  9'sd53;
	icos_lut[1874] =  9'sd128;
	qsin_lut[1875] =  9'sd77;
	icos_lut[1875] =  9'sd116;
	qsin_lut[1876] =  9'sd98;
	icos_lut[1876] =  9'sd98;
	qsin_lut[1877] =  9'sd116;
	icos_lut[1877] =  9'sd77;
	qsin_lut[1878] =  9'sd128;
	icos_lut[1878] =  9'sd53;
	qsin_lut[1879] =  9'sd136;
	icos_lut[1879] =  9'sd27;
	qsin_lut[1880] =  9'sd139;
	icos_lut[1880] =  9'sd0;
	qsin_lut[1881] =  9'sd136;
	icos_lut[1881] = -9'sd27;
	qsin_lut[1882] =  9'sd128;
	icos_lut[1882] = -9'sd53;
	qsin_lut[1883] =  9'sd116;
	icos_lut[1883] = -9'sd77;
	qsin_lut[1884] =  9'sd98;
	icos_lut[1884] = -9'sd98;
	qsin_lut[1885] =  9'sd77;
	icos_lut[1885] = -9'sd116;
	qsin_lut[1886] =  9'sd53;
	icos_lut[1886] = -9'sd128;
	qsin_lut[1887] =  9'sd27;
	icos_lut[1887] = -9'sd136;
	qsin_lut[1888] =  9'sd0;
	icos_lut[1888] = -9'sd137;
	qsin_lut[1889] = -9'sd27;
	icos_lut[1889] = -9'sd134;
	qsin_lut[1890] = -9'sd52;
	icos_lut[1890] = -9'sd127;
	qsin_lut[1891] = -9'sd76;
	icos_lut[1891] = -9'sd114;
	qsin_lut[1892] = -9'sd97;
	icos_lut[1892] = -9'sd97;
	qsin_lut[1893] = -9'sd114;
	icos_lut[1893] = -9'sd76;
	qsin_lut[1894] = -9'sd127;
	icos_lut[1894] = -9'sd52;
	qsin_lut[1895] = -9'sd134;
	icos_lut[1895] = -9'sd27;
	qsin_lut[1896] = -9'sd137;
	icos_lut[1896] = -9'sd0;
	qsin_lut[1897] = -9'sd134;
	icos_lut[1897] =  9'sd27;
	qsin_lut[1898] = -9'sd127;
	icos_lut[1898] =  9'sd52;
	qsin_lut[1899] = -9'sd114;
	icos_lut[1899] =  9'sd76;
	qsin_lut[1900] = -9'sd97;
	icos_lut[1900] =  9'sd97;
	qsin_lut[1901] = -9'sd76;
	icos_lut[1901] =  9'sd114;
	qsin_lut[1902] = -9'sd52;
	icos_lut[1902] =  9'sd127;
	qsin_lut[1903] = -9'sd27;
	icos_lut[1903] =  9'sd134;
	qsin_lut[1904] = -9'sd0;
	icos_lut[1904] =  9'sd137;
	qsin_lut[1905] =  9'sd27;
	icos_lut[1905] =  9'sd134;
	qsin_lut[1906] =  9'sd52;
	icos_lut[1906] =  9'sd127;
	qsin_lut[1907] =  9'sd76;
	icos_lut[1907] =  9'sd114;
	qsin_lut[1908] =  9'sd97;
	icos_lut[1908] =  9'sd97;
	qsin_lut[1909] =  9'sd114;
	icos_lut[1909] =  9'sd76;
	qsin_lut[1910] =  9'sd127;
	icos_lut[1910] =  9'sd52;
	qsin_lut[1911] =  9'sd134;
	icos_lut[1911] =  9'sd27;
	qsin_lut[1912] =  9'sd137;
	icos_lut[1912] =  9'sd0;
	qsin_lut[1913] =  9'sd134;
	icos_lut[1913] = -9'sd27;
	qsin_lut[1914] =  9'sd127;
	icos_lut[1914] = -9'sd52;
	qsin_lut[1915] =  9'sd114;
	icos_lut[1915] = -9'sd76;
	qsin_lut[1916] =  9'sd97;
	icos_lut[1916] = -9'sd97;
	qsin_lut[1917] =  9'sd76;
	icos_lut[1917] = -9'sd114;
	qsin_lut[1918] =  9'sd52;
	icos_lut[1918] = -9'sd127;
	qsin_lut[1919] =  9'sd27;
	icos_lut[1919] = -9'sd134;
	qsin_lut[1920] =  9'sd0;
	icos_lut[1920] = -9'sd135;
	qsin_lut[1921] = -9'sd26;
	icos_lut[1921] = -9'sd132;
	qsin_lut[1922] = -9'sd52;
	icos_lut[1922] = -9'sd125;
	qsin_lut[1923] = -9'sd75;
	icos_lut[1923] = -9'sd112;
	qsin_lut[1924] = -9'sd95;
	icos_lut[1924] = -9'sd95;
	qsin_lut[1925] = -9'sd112;
	icos_lut[1925] = -9'sd75;
	qsin_lut[1926] = -9'sd125;
	icos_lut[1926] = -9'sd52;
	qsin_lut[1927] = -9'sd132;
	icos_lut[1927] = -9'sd26;
	qsin_lut[1928] = -9'sd135;
	icos_lut[1928] = -9'sd0;
	qsin_lut[1929] = -9'sd132;
	icos_lut[1929] =  9'sd26;
	qsin_lut[1930] = -9'sd125;
	icos_lut[1930] =  9'sd52;
	qsin_lut[1931] = -9'sd112;
	icos_lut[1931] =  9'sd75;
	qsin_lut[1932] = -9'sd95;
	icos_lut[1932] =  9'sd95;
	qsin_lut[1933] = -9'sd75;
	icos_lut[1933] =  9'sd112;
	qsin_lut[1934] = -9'sd52;
	icos_lut[1934] =  9'sd125;
	qsin_lut[1935] = -9'sd26;
	icos_lut[1935] =  9'sd132;
	qsin_lut[1936] = -9'sd0;
	icos_lut[1936] =  9'sd135;
	qsin_lut[1937] =  9'sd26;
	icos_lut[1937] =  9'sd132;
	qsin_lut[1938] =  9'sd52;
	icos_lut[1938] =  9'sd125;
	qsin_lut[1939] =  9'sd75;
	icos_lut[1939] =  9'sd112;
	qsin_lut[1940] =  9'sd95;
	icos_lut[1940] =  9'sd95;
	qsin_lut[1941] =  9'sd112;
	icos_lut[1941] =  9'sd75;
	qsin_lut[1942] =  9'sd125;
	icos_lut[1942] =  9'sd52;
	qsin_lut[1943] =  9'sd132;
	icos_lut[1943] =  9'sd26;
	qsin_lut[1944] =  9'sd135;
	icos_lut[1944] =  9'sd0;
	qsin_lut[1945] =  9'sd132;
	icos_lut[1945] = -9'sd26;
	qsin_lut[1946] =  9'sd125;
	icos_lut[1946] = -9'sd52;
	qsin_lut[1947] =  9'sd112;
	icos_lut[1947] = -9'sd75;
	qsin_lut[1948] =  9'sd95;
	icos_lut[1948] = -9'sd95;
	qsin_lut[1949] =  9'sd75;
	icos_lut[1949] = -9'sd112;
	qsin_lut[1950] =  9'sd52;
	icos_lut[1950] = -9'sd125;
	qsin_lut[1951] =  9'sd26;
	icos_lut[1951] = -9'sd132;
	qsin_lut[1952] =  9'sd0;
	icos_lut[1952] = -9'sd133;
	qsin_lut[1953] = -9'sd26;
	icos_lut[1953] = -9'sd130;
	qsin_lut[1954] = -9'sd51;
	icos_lut[1954] = -9'sd123;
	qsin_lut[1955] = -9'sd74;
	icos_lut[1955] = -9'sd111;
	qsin_lut[1956] = -9'sd94;
	icos_lut[1956] = -9'sd94;
	qsin_lut[1957] = -9'sd111;
	icos_lut[1957] = -9'sd74;
	qsin_lut[1958] = -9'sd123;
	icos_lut[1958] = -9'sd51;
	qsin_lut[1959] = -9'sd130;
	icos_lut[1959] = -9'sd26;
	qsin_lut[1960] = -9'sd133;
	icos_lut[1960] = -9'sd0;
	qsin_lut[1961] = -9'sd130;
	icos_lut[1961] =  9'sd26;
	qsin_lut[1962] = -9'sd123;
	icos_lut[1962] =  9'sd51;
	qsin_lut[1963] = -9'sd111;
	icos_lut[1963] =  9'sd74;
	qsin_lut[1964] = -9'sd94;
	icos_lut[1964] =  9'sd94;
	qsin_lut[1965] = -9'sd74;
	icos_lut[1965] =  9'sd111;
	qsin_lut[1966] = -9'sd51;
	icos_lut[1966] =  9'sd123;
	qsin_lut[1967] = -9'sd26;
	icos_lut[1967] =  9'sd130;
	qsin_lut[1968] = -9'sd0;
	icos_lut[1968] =  9'sd133;
	qsin_lut[1969] =  9'sd26;
	icos_lut[1969] =  9'sd130;
	qsin_lut[1970] =  9'sd51;
	icos_lut[1970] =  9'sd123;
	qsin_lut[1971] =  9'sd74;
	icos_lut[1971] =  9'sd111;
	qsin_lut[1972] =  9'sd94;
	icos_lut[1972] =  9'sd94;
	qsin_lut[1973] =  9'sd111;
	icos_lut[1973] =  9'sd74;
	qsin_lut[1974] =  9'sd123;
	icos_lut[1974] =  9'sd51;
	qsin_lut[1975] =  9'sd130;
	icos_lut[1975] =  9'sd26;
	qsin_lut[1976] =  9'sd133;
	icos_lut[1976] =  9'sd0;
	qsin_lut[1977] =  9'sd130;
	icos_lut[1977] = -9'sd26;
	qsin_lut[1978] =  9'sd123;
	icos_lut[1978] = -9'sd51;
	qsin_lut[1979] =  9'sd111;
	icos_lut[1979] = -9'sd74;
	qsin_lut[1980] =  9'sd94;
	icos_lut[1980] = -9'sd94;
	qsin_lut[1981] =  9'sd74;
	icos_lut[1981] = -9'sd111;
	qsin_lut[1982] =  9'sd51;
	icos_lut[1982] = -9'sd123;
	qsin_lut[1983] =  9'sd26;
	icos_lut[1983] = -9'sd130;
	qsin_lut[1984] =  9'sd0;
	icos_lut[1984] = -9'sd131;
	qsin_lut[1985] = -9'sd26;
	icos_lut[1985] = -9'sd128;
	qsin_lut[1986] = -9'sd50;
	icos_lut[1986] = -9'sd121;
	qsin_lut[1987] = -9'sd73;
	icos_lut[1987] = -9'sd109;
	qsin_lut[1988] = -9'sd93;
	icos_lut[1988] = -9'sd93;
	qsin_lut[1989] = -9'sd109;
	icos_lut[1989] = -9'sd73;
	qsin_lut[1990] = -9'sd121;
	icos_lut[1990] = -9'sd50;
	qsin_lut[1991] = -9'sd128;
	icos_lut[1991] = -9'sd26;
	qsin_lut[1992] = -9'sd131;
	icos_lut[1992] = -9'sd0;
	qsin_lut[1993] = -9'sd128;
	icos_lut[1993] =  9'sd26;
	qsin_lut[1994] = -9'sd121;
	icos_lut[1994] =  9'sd50;
	qsin_lut[1995] = -9'sd109;
	icos_lut[1995] =  9'sd73;
	qsin_lut[1996] = -9'sd93;
	icos_lut[1996] =  9'sd93;
	qsin_lut[1997] = -9'sd73;
	icos_lut[1997] =  9'sd109;
	qsin_lut[1998] = -9'sd50;
	icos_lut[1998] =  9'sd121;
	qsin_lut[1999] = -9'sd26;
	icos_lut[1999] =  9'sd128;
	qsin_lut[2000] = -9'sd0;
	icos_lut[2000] =  9'sd131;
	qsin_lut[2001] =  9'sd26;
	icos_lut[2001] =  9'sd128;
	qsin_lut[2002] =  9'sd50;
	icos_lut[2002] =  9'sd121;
	qsin_lut[2003] =  9'sd73;
	icos_lut[2003] =  9'sd109;
	qsin_lut[2004] =  9'sd93;
	icos_lut[2004] =  9'sd93;
	qsin_lut[2005] =  9'sd109;
	icos_lut[2005] =  9'sd73;
	qsin_lut[2006] =  9'sd121;
	icos_lut[2006] =  9'sd50;
	qsin_lut[2007] =  9'sd128;
	icos_lut[2007] =  9'sd26;
	qsin_lut[2008] =  9'sd131;
	icos_lut[2008] =  9'sd0;
	qsin_lut[2009] =  9'sd128;
	icos_lut[2009] = -9'sd26;
	qsin_lut[2010] =  9'sd121;
	icos_lut[2010] = -9'sd50;
	qsin_lut[2011] =  9'sd109;
	icos_lut[2011] = -9'sd73;
	qsin_lut[2012] =  9'sd93;
	icos_lut[2012] = -9'sd93;
	qsin_lut[2013] =  9'sd73;
	icos_lut[2013] = -9'sd109;
	qsin_lut[2014] =  9'sd50;
	icos_lut[2014] = -9'sd121;
	qsin_lut[2015] =  9'sd26;
	icos_lut[2015] = -9'sd128;
	qsin_lut[2016] =  9'sd0;
	icos_lut[2016] = -9'sd129;
	qsin_lut[2017] = -9'sd25;
	icos_lut[2017] = -9'sd127;
	qsin_lut[2018] = -9'sd49;
	icos_lut[2018] = -9'sd119;
	qsin_lut[2019] = -9'sd72;
	icos_lut[2019] = -9'sd107;
	qsin_lut[2020] = -9'sd91;
	icos_lut[2020] = -9'sd91;
	qsin_lut[2021] = -9'sd107;
	icos_lut[2021] = -9'sd72;
	qsin_lut[2022] = -9'sd119;
	icos_lut[2022] = -9'sd49;
	qsin_lut[2023] = -9'sd127;
	icos_lut[2023] = -9'sd25;
	qsin_lut[2024] = -9'sd129;
	icos_lut[2024] = -9'sd0;
	qsin_lut[2025] = -9'sd127;
	icos_lut[2025] =  9'sd25;
	qsin_lut[2026] = -9'sd119;
	icos_lut[2026] =  9'sd49;
	qsin_lut[2027] = -9'sd107;
	icos_lut[2027] =  9'sd72;
	qsin_lut[2028] = -9'sd91;
	icos_lut[2028] =  9'sd91;
	qsin_lut[2029] = -9'sd72;
	icos_lut[2029] =  9'sd107;
	qsin_lut[2030] = -9'sd49;
	icos_lut[2030] =  9'sd119;
	qsin_lut[2031] = -9'sd25;
	icos_lut[2031] =  9'sd127;
	qsin_lut[2032] = -9'sd0;
	icos_lut[2032] =  9'sd129;
	qsin_lut[2033] =  9'sd25;
	icos_lut[2033] =  9'sd127;
	qsin_lut[2034] =  9'sd49;
	icos_lut[2034] =  9'sd119;
	qsin_lut[2035] =  9'sd72;
	icos_lut[2035] =  9'sd107;
	qsin_lut[2036] =  9'sd91;
	icos_lut[2036] =  9'sd91;
	qsin_lut[2037] =  9'sd107;
	icos_lut[2037] =  9'sd72;
	qsin_lut[2038] =  9'sd119;
	icos_lut[2038] =  9'sd49;
	qsin_lut[2039] =  9'sd127;
	icos_lut[2039] =  9'sd25;
	qsin_lut[2040] =  9'sd129;
	icos_lut[2040] =  9'sd0;
	qsin_lut[2041] =  9'sd127;
	icos_lut[2041] = -9'sd25;
	qsin_lut[2042] =  9'sd119;
	icos_lut[2042] = -9'sd49;
	qsin_lut[2043] =  9'sd107;
	icos_lut[2043] = -9'sd72;
	qsin_lut[2044] =  9'sd91;
	icos_lut[2044] = -9'sd91;
	qsin_lut[2045] =  9'sd72;
	icos_lut[2045] = -9'sd107;
	qsin_lut[2046] =  9'sd49;
	icos_lut[2046] = -9'sd119;
	qsin_lut[2047] =  9'sd25;
	icos_lut[2047] = -9'sd127;
	qsin_lut[2048] =  9'sd0;
	icos_lut[2048] = -9'sd127;
	qsin_lut[2049] = -9'sd25;
	icos_lut[2049] = -9'sd125;
	qsin_lut[2050] = -9'sd49;
	icos_lut[2050] = -9'sd117;
	qsin_lut[2051] = -9'sd71;
	icos_lut[2051] = -9'sd106;
	qsin_lut[2052] = -9'sd90;
	icos_lut[2052] = -9'sd90;
	qsin_lut[2053] = -9'sd106;
	icos_lut[2053] = -9'sd71;
	qsin_lut[2054] = -9'sd117;
	icos_lut[2054] = -9'sd49;
	qsin_lut[2055] = -9'sd125;
	icos_lut[2055] = -9'sd25;
	qsin_lut[2056] = -9'sd127;
	icos_lut[2056] = -9'sd0;
	qsin_lut[2057] = -9'sd125;
	icos_lut[2057] =  9'sd25;
	qsin_lut[2058] = -9'sd117;
	icos_lut[2058] =  9'sd49;
	qsin_lut[2059] = -9'sd106;
	icos_lut[2059] =  9'sd71;
	qsin_lut[2060] = -9'sd90;
	icos_lut[2060] =  9'sd90;
	qsin_lut[2061] = -9'sd71;
	icos_lut[2061] =  9'sd106;
	qsin_lut[2062] = -9'sd49;
	icos_lut[2062] =  9'sd117;
	qsin_lut[2063] = -9'sd25;
	icos_lut[2063] =  9'sd125;
	qsin_lut[2064] = -9'sd0;
	icos_lut[2064] =  9'sd127;
	qsin_lut[2065] =  9'sd25;
	icos_lut[2065] =  9'sd125;
	qsin_lut[2066] =  9'sd49;
	icos_lut[2066] =  9'sd117;
	qsin_lut[2067] =  9'sd71;
	icos_lut[2067] =  9'sd106;
	qsin_lut[2068] =  9'sd90;
	icos_lut[2068] =  9'sd90;
	qsin_lut[2069] =  9'sd106;
	icos_lut[2069] =  9'sd71;
	qsin_lut[2070] =  9'sd117;
	icos_lut[2070] =  9'sd49;
	qsin_lut[2071] =  9'sd125;
	icos_lut[2071] =  9'sd25;
	qsin_lut[2072] =  9'sd127;
	icos_lut[2072] =  9'sd0;
	qsin_lut[2073] =  9'sd125;
	icos_lut[2073] = -9'sd25;
	qsin_lut[2074] =  9'sd117;
	icos_lut[2074] = -9'sd49;
	qsin_lut[2075] =  9'sd106;
	icos_lut[2075] = -9'sd71;
	qsin_lut[2076] =  9'sd90;
	icos_lut[2076] = -9'sd90;
	qsin_lut[2077] =  9'sd71;
	icos_lut[2077] = -9'sd106;
	qsin_lut[2078] =  9'sd49;
	icos_lut[2078] = -9'sd117;
	qsin_lut[2079] =  9'sd25;
	icos_lut[2079] = -9'sd125;
	qsin_lut[2080] =  9'sd0;
	icos_lut[2080] = -9'sd125;
	qsin_lut[2081] = -9'sd24;
	icos_lut[2081] = -9'sd123;
	qsin_lut[2082] = -9'sd48;
	icos_lut[2082] = -9'sd115;
	qsin_lut[2083] = -9'sd69;
	icos_lut[2083] = -9'sd104;
	qsin_lut[2084] = -9'sd88;
	icos_lut[2084] = -9'sd88;
	qsin_lut[2085] = -9'sd104;
	icos_lut[2085] = -9'sd69;
	qsin_lut[2086] = -9'sd115;
	icos_lut[2086] = -9'sd48;
	qsin_lut[2087] = -9'sd123;
	icos_lut[2087] = -9'sd24;
	qsin_lut[2088] = -9'sd125;
	icos_lut[2088] = -9'sd0;
	qsin_lut[2089] = -9'sd123;
	icos_lut[2089] =  9'sd24;
	qsin_lut[2090] = -9'sd115;
	icos_lut[2090] =  9'sd48;
	qsin_lut[2091] = -9'sd104;
	icos_lut[2091] =  9'sd69;
	qsin_lut[2092] = -9'sd88;
	icos_lut[2092] =  9'sd88;
	qsin_lut[2093] = -9'sd69;
	icos_lut[2093] =  9'sd104;
	qsin_lut[2094] = -9'sd48;
	icos_lut[2094] =  9'sd115;
	qsin_lut[2095] = -9'sd24;
	icos_lut[2095] =  9'sd123;
	qsin_lut[2096] = -9'sd0;
	icos_lut[2096] =  9'sd125;
	qsin_lut[2097] =  9'sd24;
	icos_lut[2097] =  9'sd123;
	qsin_lut[2098] =  9'sd48;
	icos_lut[2098] =  9'sd115;
	qsin_lut[2099] =  9'sd69;
	icos_lut[2099] =  9'sd104;
	qsin_lut[2100] =  9'sd88;
	icos_lut[2100] =  9'sd88;
	qsin_lut[2101] =  9'sd104;
	icos_lut[2101] =  9'sd69;
	qsin_lut[2102] =  9'sd115;
	icos_lut[2102] =  9'sd48;
	qsin_lut[2103] =  9'sd123;
	icos_lut[2103] =  9'sd24;
	qsin_lut[2104] =  9'sd125;
	icos_lut[2104] =  9'sd0;
	qsin_lut[2105] =  9'sd123;
	icos_lut[2105] = -9'sd24;
	qsin_lut[2106] =  9'sd115;
	icos_lut[2106] = -9'sd48;
	qsin_lut[2107] =  9'sd104;
	icos_lut[2107] = -9'sd69;
	qsin_lut[2108] =  9'sd88;
	icos_lut[2108] = -9'sd88;
	qsin_lut[2109] =  9'sd69;
	icos_lut[2109] = -9'sd104;
	qsin_lut[2110] =  9'sd48;
	icos_lut[2110] = -9'sd115;
	qsin_lut[2111] =  9'sd24;
	icos_lut[2111] = -9'sd123;
	qsin_lut[2112] =  9'sd0;
	icos_lut[2112] = -9'sd123;
	qsin_lut[2113] = -9'sd24;
	icos_lut[2113] = -9'sd121;
	qsin_lut[2114] = -9'sd47;
	icos_lut[2114] = -9'sd114;
	qsin_lut[2115] = -9'sd68;
	icos_lut[2115] = -9'sd102;
	qsin_lut[2116] = -9'sd87;
	icos_lut[2116] = -9'sd87;
	qsin_lut[2117] = -9'sd102;
	icos_lut[2117] = -9'sd68;
	qsin_lut[2118] = -9'sd114;
	icos_lut[2118] = -9'sd47;
	qsin_lut[2119] = -9'sd121;
	icos_lut[2119] = -9'sd24;
	qsin_lut[2120] = -9'sd123;
	icos_lut[2120] = -9'sd0;
	qsin_lut[2121] = -9'sd121;
	icos_lut[2121] =  9'sd24;
	qsin_lut[2122] = -9'sd114;
	icos_lut[2122] =  9'sd47;
	qsin_lut[2123] = -9'sd102;
	icos_lut[2123] =  9'sd68;
	qsin_lut[2124] = -9'sd87;
	icos_lut[2124] =  9'sd87;
	qsin_lut[2125] = -9'sd68;
	icos_lut[2125] =  9'sd102;
	qsin_lut[2126] = -9'sd47;
	icos_lut[2126] =  9'sd114;
	qsin_lut[2127] = -9'sd24;
	icos_lut[2127] =  9'sd121;
	qsin_lut[2128] = -9'sd0;
	icos_lut[2128] =  9'sd123;
	qsin_lut[2129] =  9'sd24;
	icos_lut[2129] =  9'sd121;
	qsin_lut[2130] =  9'sd47;
	icos_lut[2130] =  9'sd114;
	qsin_lut[2131] =  9'sd68;
	icos_lut[2131] =  9'sd102;
	qsin_lut[2132] =  9'sd87;
	icos_lut[2132] =  9'sd87;
	qsin_lut[2133] =  9'sd102;
	icos_lut[2133] =  9'sd68;
	qsin_lut[2134] =  9'sd114;
	icos_lut[2134] =  9'sd47;
	qsin_lut[2135] =  9'sd121;
	icos_lut[2135] =  9'sd24;
	qsin_lut[2136] =  9'sd123;
	icos_lut[2136] =  9'sd0;
	qsin_lut[2137] =  9'sd121;
	icos_lut[2137] = -9'sd24;
	qsin_lut[2138] =  9'sd114;
	icos_lut[2138] = -9'sd47;
	qsin_lut[2139] =  9'sd102;
	icos_lut[2139] = -9'sd68;
	qsin_lut[2140] =  9'sd87;
	icos_lut[2140] = -9'sd87;
	qsin_lut[2141] =  9'sd68;
	icos_lut[2141] = -9'sd102;
	qsin_lut[2142] =  9'sd47;
	icos_lut[2142] = -9'sd114;
	qsin_lut[2143] =  9'sd24;
	icos_lut[2143] = -9'sd121;
	qsin_lut[2144] =  9'sd0;
	icos_lut[2144] = -9'sd121;
	qsin_lut[2145] = -9'sd24;
	icos_lut[2145] = -9'sd119;
	qsin_lut[2146] = -9'sd46;
	icos_lut[2146] = -9'sd112;
	qsin_lut[2147] = -9'sd67;
	icos_lut[2147] = -9'sd101;
	qsin_lut[2148] = -9'sd86;
	icos_lut[2148] = -9'sd86;
	qsin_lut[2149] = -9'sd101;
	icos_lut[2149] = -9'sd67;
	qsin_lut[2150] = -9'sd112;
	icos_lut[2150] = -9'sd46;
	qsin_lut[2151] = -9'sd119;
	icos_lut[2151] = -9'sd24;
	qsin_lut[2152] = -9'sd121;
	icos_lut[2152] = -9'sd0;
	qsin_lut[2153] = -9'sd119;
	icos_lut[2153] =  9'sd24;
	qsin_lut[2154] = -9'sd112;
	icos_lut[2154] =  9'sd46;
	qsin_lut[2155] = -9'sd101;
	icos_lut[2155] =  9'sd67;
	qsin_lut[2156] = -9'sd86;
	icos_lut[2156] =  9'sd86;
	qsin_lut[2157] = -9'sd67;
	icos_lut[2157] =  9'sd101;
	qsin_lut[2158] = -9'sd46;
	icos_lut[2158] =  9'sd112;
	qsin_lut[2159] = -9'sd24;
	icos_lut[2159] =  9'sd119;
	qsin_lut[2160] = -9'sd0;
	icos_lut[2160] =  9'sd121;
	qsin_lut[2161] =  9'sd24;
	icos_lut[2161] =  9'sd119;
	qsin_lut[2162] =  9'sd46;
	icos_lut[2162] =  9'sd112;
	qsin_lut[2163] =  9'sd67;
	icos_lut[2163] =  9'sd101;
	qsin_lut[2164] =  9'sd86;
	icos_lut[2164] =  9'sd86;
	qsin_lut[2165] =  9'sd101;
	icos_lut[2165] =  9'sd67;
	qsin_lut[2166] =  9'sd112;
	icos_lut[2166] =  9'sd46;
	qsin_lut[2167] =  9'sd119;
	icos_lut[2167] =  9'sd24;
	qsin_lut[2168] =  9'sd121;
	icos_lut[2168] =  9'sd0;
	qsin_lut[2169] =  9'sd119;
	icos_lut[2169] = -9'sd24;
	qsin_lut[2170] =  9'sd112;
	icos_lut[2170] = -9'sd46;
	qsin_lut[2171] =  9'sd101;
	icos_lut[2171] = -9'sd67;
	qsin_lut[2172] =  9'sd86;
	icos_lut[2172] = -9'sd86;
	qsin_lut[2173] =  9'sd67;
	icos_lut[2173] = -9'sd101;
	qsin_lut[2174] =  9'sd46;
	icos_lut[2174] = -9'sd112;
	qsin_lut[2175] =  9'sd24;
	icos_lut[2175] = -9'sd119;
	qsin_lut[2176] =  9'sd0;
	icos_lut[2176] = -9'sd119;
	qsin_lut[2177] = -9'sd23;
	icos_lut[2177] = -9'sd117;
	qsin_lut[2178] = -9'sd46;
	icos_lut[2178] = -9'sd110;
	qsin_lut[2179] = -9'sd66;
	icos_lut[2179] = -9'sd99;
	qsin_lut[2180] = -9'sd84;
	icos_lut[2180] = -9'sd84;
	qsin_lut[2181] = -9'sd99;
	icos_lut[2181] = -9'sd66;
	qsin_lut[2182] = -9'sd110;
	icos_lut[2182] = -9'sd46;
	qsin_lut[2183] = -9'sd117;
	icos_lut[2183] = -9'sd23;
	qsin_lut[2184] = -9'sd119;
	icos_lut[2184] = -9'sd0;
	qsin_lut[2185] = -9'sd117;
	icos_lut[2185] =  9'sd23;
	qsin_lut[2186] = -9'sd110;
	icos_lut[2186] =  9'sd46;
	qsin_lut[2187] = -9'sd99;
	icos_lut[2187] =  9'sd66;
	qsin_lut[2188] = -9'sd84;
	icos_lut[2188] =  9'sd84;
	qsin_lut[2189] = -9'sd66;
	icos_lut[2189] =  9'sd99;
	qsin_lut[2190] = -9'sd46;
	icos_lut[2190] =  9'sd110;
	qsin_lut[2191] = -9'sd23;
	icos_lut[2191] =  9'sd117;
	qsin_lut[2192] = -9'sd0;
	icos_lut[2192] =  9'sd119;
	qsin_lut[2193] =  9'sd23;
	icos_lut[2193] =  9'sd117;
	qsin_lut[2194] =  9'sd46;
	icos_lut[2194] =  9'sd110;
	qsin_lut[2195] =  9'sd66;
	icos_lut[2195] =  9'sd99;
	qsin_lut[2196] =  9'sd84;
	icos_lut[2196] =  9'sd84;
	qsin_lut[2197] =  9'sd99;
	icos_lut[2197] =  9'sd66;
	qsin_lut[2198] =  9'sd110;
	icos_lut[2198] =  9'sd46;
	qsin_lut[2199] =  9'sd117;
	icos_lut[2199] =  9'sd23;
	qsin_lut[2200] =  9'sd119;
	icos_lut[2200] =  9'sd0;
	qsin_lut[2201] =  9'sd117;
	icos_lut[2201] = -9'sd23;
	qsin_lut[2202] =  9'sd110;
	icos_lut[2202] = -9'sd46;
	qsin_lut[2203] =  9'sd99;
	icos_lut[2203] = -9'sd66;
	qsin_lut[2204] =  9'sd84;
	icos_lut[2204] = -9'sd84;
	qsin_lut[2205] =  9'sd66;
	icos_lut[2205] = -9'sd99;
	qsin_lut[2206] =  9'sd46;
	icos_lut[2206] = -9'sd110;
	qsin_lut[2207] =  9'sd23;
	icos_lut[2207] = -9'sd117;
	qsin_lut[2208] =  9'sd0;
	icos_lut[2208] = -9'sd117;
	qsin_lut[2209] = -9'sd23;
	icos_lut[2209] = -9'sd115;
	qsin_lut[2210] = -9'sd45;
	icos_lut[2210] = -9'sd108;
	qsin_lut[2211] = -9'sd65;
	icos_lut[2211] = -9'sd97;
	qsin_lut[2212] = -9'sd83;
	icos_lut[2212] = -9'sd83;
	qsin_lut[2213] = -9'sd97;
	icos_lut[2213] = -9'sd65;
	qsin_lut[2214] = -9'sd108;
	icos_lut[2214] = -9'sd45;
	qsin_lut[2215] = -9'sd115;
	icos_lut[2215] = -9'sd23;
	qsin_lut[2216] = -9'sd117;
	icos_lut[2216] = -9'sd0;
	qsin_lut[2217] = -9'sd115;
	icos_lut[2217] =  9'sd23;
	qsin_lut[2218] = -9'sd108;
	icos_lut[2218] =  9'sd45;
	qsin_lut[2219] = -9'sd97;
	icos_lut[2219] =  9'sd65;
	qsin_lut[2220] = -9'sd83;
	icos_lut[2220] =  9'sd83;
	qsin_lut[2221] = -9'sd65;
	icos_lut[2221] =  9'sd97;
	qsin_lut[2222] = -9'sd45;
	icos_lut[2222] =  9'sd108;
	qsin_lut[2223] = -9'sd23;
	icos_lut[2223] =  9'sd115;
	qsin_lut[2224] = -9'sd0;
	icos_lut[2224] =  9'sd117;
	qsin_lut[2225] =  9'sd23;
	icos_lut[2225] =  9'sd115;
	qsin_lut[2226] =  9'sd45;
	icos_lut[2226] =  9'sd108;
	qsin_lut[2227] =  9'sd65;
	icos_lut[2227] =  9'sd97;
	qsin_lut[2228] =  9'sd83;
	icos_lut[2228] =  9'sd83;
	qsin_lut[2229] =  9'sd97;
	icos_lut[2229] =  9'sd65;
	qsin_lut[2230] =  9'sd108;
	icos_lut[2230] =  9'sd45;
	qsin_lut[2231] =  9'sd115;
	icos_lut[2231] =  9'sd23;
	qsin_lut[2232] =  9'sd117;
	icos_lut[2232] =  9'sd0;
	qsin_lut[2233] =  9'sd115;
	icos_lut[2233] = -9'sd23;
	qsin_lut[2234] =  9'sd108;
	icos_lut[2234] = -9'sd45;
	qsin_lut[2235] =  9'sd97;
	icos_lut[2235] = -9'sd65;
	qsin_lut[2236] =  9'sd83;
	icos_lut[2236] = -9'sd83;
	qsin_lut[2237] =  9'sd65;
	icos_lut[2237] = -9'sd97;
	qsin_lut[2238] =  9'sd45;
	icos_lut[2238] = -9'sd108;
	qsin_lut[2239] =  9'sd23;
	icos_lut[2239] = -9'sd115;
	qsin_lut[2240] =  9'sd0;
	icos_lut[2240] = -9'sd115;
	qsin_lut[2241] = -9'sd22;
	icos_lut[2241] = -9'sd113;
	qsin_lut[2242] = -9'sd44;
	icos_lut[2242] = -9'sd106;
	qsin_lut[2243] = -9'sd64;
	icos_lut[2243] = -9'sd96;
	qsin_lut[2244] = -9'sd81;
	icos_lut[2244] = -9'sd81;
	qsin_lut[2245] = -9'sd96;
	icos_lut[2245] = -9'sd64;
	qsin_lut[2246] = -9'sd106;
	icos_lut[2246] = -9'sd44;
	qsin_lut[2247] = -9'sd113;
	icos_lut[2247] = -9'sd22;
	qsin_lut[2248] = -9'sd115;
	icos_lut[2248] = -9'sd0;
	qsin_lut[2249] = -9'sd113;
	icos_lut[2249] =  9'sd22;
	qsin_lut[2250] = -9'sd106;
	icos_lut[2250] =  9'sd44;
	qsin_lut[2251] = -9'sd96;
	icos_lut[2251] =  9'sd64;
	qsin_lut[2252] = -9'sd81;
	icos_lut[2252] =  9'sd81;
	qsin_lut[2253] = -9'sd64;
	icos_lut[2253] =  9'sd96;
	qsin_lut[2254] = -9'sd44;
	icos_lut[2254] =  9'sd106;
	qsin_lut[2255] = -9'sd22;
	icos_lut[2255] =  9'sd113;
	qsin_lut[2256] = -9'sd0;
	icos_lut[2256] =  9'sd115;
	qsin_lut[2257] =  9'sd22;
	icos_lut[2257] =  9'sd113;
	qsin_lut[2258] =  9'sd44;
	icos_lut[2258] =  9'sd106;
	qsin_lut[2259] =  9'sd64;
	icos_lut[2259] =  9'sd96;
	qsin_lut[2260] =  9'sd81;
	icos_lut[2260] =  9'sd81;
	qsin_lut[2261] =  9'sd96;
	icos_lut[2261] =  9'sd64;
	qsin_lut[2262] =  9'sd106;
	icos_lut[2262] =  9'sd44;
	qsin_lut[2263] =  9'sd113;
	icos_lut[2263] =  9'sd22;
	qsin_lut[2264] =  9'sd115;
	icos_lut[2264] =  9'sd0;
	qsin_lut[2265] =  9'sd113;
	icos_lut[2265] = -9'sd22;
	qsin_lut[2266] =  9'sd106;
	icos_lut[2266] = -9'sd44;
	qsin_lut[2267] =  9'sd96;
	icos_lut[2267] = -9'sd64;
	qsin_lut[2268] =  9'sd81;
	icos_lut[2268] = -9'sd81;
	qsin_lut[2269] =  9'sd64;
	icos_lut[2269] = -9'sd96;
	qsin_lut[2270] =  9'sd44;
	icos_lut[2270] = -9'sd106;
	qsin_lut[2271] =  9'sd22;
	icos_lut[2271] = -9'sd113;
	qsin_lut[2272] =  9'sd0;
	icos_lut[2272] = -9'sd113;
	qsin_lut[2273] = -9'sd22;
	icos_lut[2273] = -9'sd111;
	qsin_lut[2274] = -9'sd43;
	icos_lut[2274] = -9'sd104;
	qsin_lut[2275] = -9'sd63;
	icos_lut[2275] = -9'sd94;
	qsin_lut[2276] = -9'sd80;
	icos_lut[2276] = -9'sd80;
	qsin_lut[2277] = -9'sd94;
	icos_lut[2277] = -9'sd63;
	qsin_lut[2278] = -9'sd104;
	icos_lut[2278] = -9'sd43;
	qsin_lut[2279] = -9'sd111;
	icos_lut[2279] = -9'sd22;
	qsin_lut[2280] = -9'sd113;
	icos_lut[2280] = -9'sd0;
	qsin_lut[2281] = -9'sd111;
	icos_lut[2281] =  9'sd22;
	qsin_lut[2282] = -9'sd104;
	icos_lut[2282] =  9'sd43;
	qsin_lut[2283] = -9'sd94;
	icos_lut[2283] =  9'sd63;
	qsin_lut[2284] = -9'sd80;
	icos_lut[2284] =  9'sd80;
	qsin_lut[2285] = -9'sd63;
	icos_lut[2285] =  9'sd94;
	qsin_lut[2286] = -9'sd43;
	icos_lut[2286] =  9'sd104;
	qsin_lut[2287] = -9'sd22;
	icos_lut[2287] =  9'sd111;
	qsin_lut[2288] = -9'sd0;
	icos_lut[2288] =  9'sd113;
	qsin_lut[2289] =  9'sd22;
	icos_lut[2289] =  9'sd111;
	qsin_lut[2290] =  9'sd43;
	icos_lut[2290] =  9'sd104;
	qsin_lut[2291] =  9'sd63;
	icos_lut[2291] =  9'sd94;
	qsin_lut[2292] =  9'sd80;
	icos_lut[2292] =  9'sd80;
	qsin_lut[2293] =  9'sd94;
	icos_lut[2293] =  9'sd63;
	qsin_lut[2294] =  9'sd104;
	icos_lut[2294] =  9'sd43;
	qsin_lut[2295] =  9'sd111;
	icos_lut[2295] =  9'sd22;
	qsin_lut[2296] =  9'sd113;
	icos_lut[2296] =  9'sd0;
	qsin_lut[2297] =  9'sd111;
	icos_lut[2297] = -9'sd22;
	qsin_lut[2298] =  9'sd104;
	icos_lut[2298] = -9'sd43;
	qsin_lut[2299] =  9'sd94;
	icos_lut[2299] = -9'sd63;
	qsin_lut[2300] =  9'sd80;
	icos_lut[2300] = -9'sd80;
	qsin_lut[2301] =  9'sd63;
	icos_lut[2301] = -9'sd94;
	qsin_lut[2302] =  9'sd43;
	icos_lut[2302] = -9'sd104;
	qsin_lut[2303] =  9'sd22;
	icos_lut[2303] = -9'sd111;
	qsin_lut[2304] =  9'sd0;
	icos_lut[2304] = -9'sd111;
	qsin_lut[2305] = -9'sd22;
	icos_lut[2305] = -9'sd109;
	qsin_lut[2306] = -9'sd42;
	icos_lut[2306] = -9'sd103;
	qsin_lut[2307] = -9'sd62;
	icos_lut[2307] = -9'sd92;
	qsin_lut[2308] = -9'sd78;
	icos_lut[2308] = -9'sd78;
	qsin_lut[2309] = -9'sd92;
	icos_lut[2309] = -9'sd62;
	qsin_lut[2310] = -9'sd103;
	icos_lut[2310] = -9'sd42;
	qsin_lut[2311] = -9'sd109;
	icos_lut[2311] = -9'sd22;
	qsin_lut[2312] = -9'sd111;
	icos_lut[2312] = -9'sd0;
	qsin_lut[2313] = -9'sd109;
	icos_lut[2313] =  9'sd22;
	qsin_lut[2314] = -9'sd103;
	icos_lut[2314] =  9'sd42;
	qsin_lut[2315] = -9'sd92;
	icos_lut[2315] =  9'sd62;
	qsin_lut[2316] = -9'sd78;
	icos_lut[2316] =  9'sd78;
	qsin_lut[2317] = -9'sd62;
	icos_lut[2317] =  9'sd92;
	qsin_lut[2318] = -9'sd42;
	icos_lut[2318] =  9'sd103;
	qsin_lut[2319] = -9'sd22;
	icos_lut[2319] =  9'sd109;
	qsin_lut[2320] = -9'sd0;
	icos_lut[2320] =  9'sd111;
	qsin_lut[2321] =  9'sd22;
	icos_lut[2321] =  9'sd109;
	qsin_lut[2322] =  9'sd42;
	icos_lut[2322] =  9'sd103;
	qsin_lut[2323] =  9'sd62;
	icos_lut[2323] =  9'sd92;
	qsin_lut[2324] =  9'sd78;
	icos_lut[2324] =  9'sd78;
	qsin_lut[2325] =  9'sd92;
	icos_lut[2325] =  9'sd62;
	qsin_lut[2326] =  9'sd103;
	icos_lut[2326] =  9'sd42;
	qsin_lut[2327] =  9'sd109;
	icos_lut[2327] =  9'sd22;
	qsin_lut[2328] =  9'sd111;
	icos_lut[2328] =  9'sd0;
	qsin_lut[2329] =  9'sd109;
	icos_lut[2329] = -9'sd22;
	qsin_lut[2330] =  9'sd103;
	icos_lut[2330] = -9'sd42;
	qsin_lut[2331] =  9'sd92;
	icos_lut[2331] = -9'sd62;
	qsin_lut[2332] =  9'sd78;
	icos_lut[2332] = -9'sd78;
	qsin_lut[2333] =  9'sd62;
	icos_lut[2333] = -9'sd92;
	qsin_lut[2334] =  9'sd42;
	icos_lut[2334] = -9'sd103;
	qsin_lut[2335] =  9'sd22;
	icos_lut[2335] = -9'sd109;
	qsin_lut[2336] =  9'sd0;
	icos_lut[2336] = -9'sd109;
	qsin_lut[2337] = -9'sd21;
	icos_lut[2337] = -9'sd107;
	qsin_lut[2338] = -9'sd42;
	icos_lut[2338] = -9'sd101;
	qsin_lut[2339] = -9'sd61;
	icos_lut[2339] = -9'sd91;
	qsin_lut[2340] = -9'sd77;
	icos_lut[2340] = -9'sd77;
	qsin_lut[2341] = -9'sd91;
	icos_lut[2341] = -9'sd61;
	qsin_lut[2342] = -9'sd101;
	icos_lut[2342] = -9'sd42;
	qsin_lut[2343] = -9'sd107;
	icos_lut[2343] = -9'sd21;
	qsin_lut[2344] = -9'sd109;
	icos_lut[2344] = -9'sd0;
	qsin_lut[2345] = -9'sd107;
	icos_lut[2345] =  9'sd21;
	qsin_lut[2346] = -9'sd101;
	icos_lut[2346] =  9'sd42;
	qsin_lut[2347] = -9'sd91;
	icos_lut[2347] =  9'sd61;
	qsin_lut[2348] = -9'sd77;
	icos_lut[2348] =  9'sd77;
	qsin_lut[2349] = -9'sd61;
	icos_lut[2349] =  9'sd91;
	qsin_lut[2350] = -9'sd42;
	icos_lut[2350] =  9'sd101;
	qsin_lut[2351] = -9'sd21;
	icos_lut[2351] =  9'sd107;
	qsin_lut[2352] = -9'sd0;
	icos_lut[2352] =  9'sd109;
	qsin_lut[2353] =  9'sd21;
	icos_lut[2353] =  9'sd107;
	qsin_lut[2354] =  9'sd42;
	icos_lut[2354] =  9'sd101;
	qsin_lut[2355] =  9'sd61;
	icos_lut[2355] =  9'sd91;
	qsin_lut[2356] =  9'sd77;
	icos_lut[2356] =  9'sd77;
	qsin_lut[2357] =  9'sd91;
	icos_lut[2357] =  9'sd61;
	qsin_lut[2358] =  9'sd101;
	icos_lut[2358] =  9'sd42;
	qsin_lut[2359] =  9'sd107;
	icos_lut[2359] =  9'sd21;
	qsin_lut[2360] =  9'sd109;
	icos_lut[2360] =  9'sd0;
	qsin_lut[2361] =  9'sd107;
	icos_lut[2361] = -9'sd21;
	qsin_lut[2362] =  9'sd101;
	icos_lut[2362] = -9'sd42;
	qsin_lut[2363] =  9'sd91;
	icos_lut[2363] = -9'sd61;
	qsin_lut[2364] =  9'sd77;
	icos_lut[2364] = -9'sd77;
	qsin_lut[2365] =  9'sd61;
	icos_lut[2365] = -9'sd91;
	qsin_lut[2366] =  9'sd42;
	icos_lut[2366] = -9'sd101;
	qsin_lut[2367] =  9'sd21;
	icos_lut[2367] = -9'sd107;
	qsin_lut[2368] =  9'sd0;
	icos_lut[2368] = -9'sd107;
	qsin_lut[2369] = -9'sd21;
	icos_lut[2369] = -9'sd105;
	qsin_lut[2370] = -9'sd41;
	icos_lut[2370] = -9'sd99;
	qsin_lut[2371] = -9'sd59;
	icos_lut[2371] = -9'sd89;
	qsin_lut[2372] = -9'sd76;
	icos_lut[2372] = -9'sd76;
	qsin_lut[2373] = -9'sd89;
	icos_lut[2373] = -9'sd59;
	qsin_lut[2374] = -9'sd99;
	icos_lut[2374] = -9'sd41;
	qsin_lut[2375] = -9'sd105;
	icos_lut[2375] = -9'sd21;
	qsin_lut[2376] = -9'sd107;
	icos_lut[2376] = -9'sd0;
	qsin_lut[2377] = -9'sd105;
	icos_lut[2377] =  9'sd21;
	qsin_lut[2378] = -9'sd99;
	icos_lut[2378] =  9'sd41;
	qsin_lut[2379] = -9'sd89;
	icos_lut[2379] =  9'sd59;
	qsin_lut[2380] = -9'sd76;
	icos_lut[2380] =  9'sd76;
	qsin_lut[2381] = -9'sd59;
	icos_lut[2381] =  9'sd89;
	qsin_lut[2382] = -9'sd41;
	icos_lut[2382] =  9'sd99;
	qsin_lut[2383] = -9'sd21;
	icos_lut[2383] =  9'sd105;
	qsin_lut[2384] = -9'sd0;
	icos_lut[2384] =  9'sd107;
	qsin_lut[2385] =  9'sd21;
	icos_lut[2385] =  9'sd105;
	qsin_lut[2386] =  9'sd41;
	icos_lut[2386] =  9'sd99;
	qsin_lut[2387] =  9'sd59;
	icos_lut[2387] =  9'sd89;
	qsin_lut[2388] =  9'sd76;
	icos_lut[2388] =  9'sd76;
	qsin_lut[2389] =  9'sd89;
	icos_lut[2389] =  9'sd59;
	qsin_lut[2390] =  9'sd99;
	icos_lut[2390] =  9'sd41;
	qsin_lut[2391] =  9'sd105;
	icos_lut[2391] =  9'sd21;
	qsin_lut[2392] =  9'sd107;
	icos_lut[2392] =  9'sd0;
	qsin_lut[2393] =  9'sd105;
	icos_lut[2393] = -9'sd21;
	qsin_lut[2394] =  9'sd99;
	icos_lut[2394] = -9'sd41;
	qsin_lut[2395] =  9'sd89;
	icos_lut[2395] = -9'sd59;
	qsin_lut[2396] =  9'sd76;
	icos_lut[2396] = -9'sd76;
	qsin_lut[2397] =  9'sd59;
	icos_lut[2397] = -9'sd89;
	qsin_lut[2398] =  9'sd41;
	icos_lut[2398] = -9'sd99;
	qsin_lut[2399] =  9'sd21;
	icos_lut[2399] = -9'sd105;
	qsin_lut[2400] =  9'sd0;
	icos_lut[2400] = -9'sd105;
	qsin_lut[2401] = -9'sd20;
	icos_lut[2401] = -9'sd103;
	qsin_lut[2402] = -9'sd40;
	icos_lut[2402] = -9'sd97;
	qsin_lut[2403] = -9'sd58;
	icos_lut[2403] = -9'sd87;
	qsin_lut[2404] = -9'sd74;
	icos_lut[2404] = -9'sd74;
	qsin_lut[2405] = -9'sd87;
	icos_lut[2405] = -9'sd58;
	qsin_lut[2406] = -9'sd97;
	icos_lut[2406] = -9'sd40;
	qsin_lut[2407] = -9'sd103;
	icos_lut[2407] = -9'sd20;
	qsin_lut[2408] = -9'sd105;
	icos_lut[2408] = -9'sd0;
	qsin_lut[2409] = -9'sd103;
	icos_lut[2409] =  9'sd20;
	qsin_lut[2410] = -9'sd97;
	icos_lut[2410] =  9'sd40;
	qsin_lut[2411] = -9'sd87;
	icos_lut[2411] =  9'sd58;
	qsin_lut[2412] = -9'sd74;
	icos_lut[2412] =  9'sd74;
	qsin_lut[2413] = -9'sd58;
	icos_lut[2413] =  9'sd87;
	qsin_lut[2414] = -9'sd40;
	icos_lut[2414] =  9'sd97;
	qsin_lut[2415] = -9'sd20;
	icos_lut[2415] =  9'sd103;
	qsin_lut[2416] = -9'sd0;
	icos_lut[2416] =  9'sd105;
	qsin_lut[2417] =  9'sd20;
	icos_lut[2417] =  9'sd103;
	qsin_lut[2418] =  9'sd40;
	icos_lut[2418] =  9'sd97;
	qsin_lut[2419] =  9'sd58;
	icos_lut[2419] =  9'sd87;
	qsin_lut[2420] =  9'sd74;
	icos_lut[2420] =  9'sd74;
	qsin_lut[2421] =  9'sd87;
	icos_lut[2421] =  9'sd58;
	qsin_lut[2422] =  9'sd97;
	icos_lut[2422] =  9'sd40;
	qsin_lut[2423] =  9'sd103;
	icos_lut[2423] =  9'sd20;
	qsin_lut[2424] =  9'sd105;
	icos_lut[2424] =  9'sd0;
	qsin_lut[2425] =  9'sd103;
	icos_lut[2425] = -9'sd20;
	qsin_lut[2426] =  9'sd97;
	icos_lut[2426] = -9'sd40;
	qsin_lut[2427] =  9'sd87;
	icos_lut[2427] = -9'sd58;
	qsin_lut[2428] =  9'sd74;
	icos_lut[2428] = -9'sd74;
	qsin_lut[2429] =  9'sd58;
	icos_lut[2429] = -9'sd87;
	qsin_lut[2430] =  9'sd40;
	icos_lut[2430] = -9'sd97;
	qsin_lut[2431] =  9'sd20;
	icos_lut[2431] = -9'sd103;
	qsin_lut[2432] =  9'sd0;
	icos_lut[2432] = -9'sd103;
	qsin_lut[2433] = -9'sd20;
	icos_lut[2433] = -9'sd101;
	qsin_lut[2434] = -9'sd39;
	icos_lut[2434] = -9'sd95;
	qsin_lut[2435] = -9'sd57;
	icos_lut[2435] = -9'sd86;
	qsin_lut[2436] = -9'sd73;
	icos_lut[2436] = -9'sd73;
	qsin_lut[2437] = -9'sd86;
	icos_lut[2437] = -9'sd57;
	qsin_lut[2438] = -9'sd95;
	icos_lut[2438] = -9'sd39;
	qsin_lut[2439] = -9'sd101;
	icos_lut[2439] = -9'sd20;
	qsin_lut[2440] = -9'sd103;
	icos_lut[2440] = -9'sd0;
	qsin_lut[2441] = -9'sd101;
	icos_lut[2441] =  9'sd20;
	qsin_lut[2442] = -9'sd95;
	icos_lut[2442] =  9'sd39;
	qsin_lut[2443] = -9'sd86;
	icos_lut[2443] =  9'sd57;
	qsin_lut[2444] = -9'sd73;
	icos_lut[2444] =  9'sd73;
	qsin_lut[2445] = -9'sd57;
	icos_lut[2445] =  9'sd86;
	qsin_lut[2446] = -9'sd39;
	icos_lut[2446] =  9'sd95;
	qsin_lut[2447] = -9'sd20;
	icos_lut[2447] =  9'sd101;
	qsin_lut[2448] = -9'sd0;
	icos_lut[2448] =  9'sd103;
	qsin_lut[2449] =  9'sd20;
	icos_lut[2449] =  9'sd101;
	qsin_lut[2450] =  9'sd39;
	icos_lut[2450] =  9'sd95;
	qsin_lut[2451] =  9'sd57;
	icos_lut[2451] =  9'sd86;
	qsin_lut[2452] =  9'sd73;
	icos_lut[2452] =  9'sd73;
	qsin_lut[2453] =  9'sd86;
	icos_lut[2453] =  9'sd57;
	qsin_lut[2454] =  9'sd95;
	icos_lut[2454] =  9'sd39;
	qsin_lut[2455] =  9'sd101;
	icos_lut[2455] =  9'sd20;
	qsin_lut[2456] =  9'sd103;
	icos_lut[2456] =  9'sd0;
	qsin_lut[2457] =  9'sd101;
	icos_lut[2457] = -9'sd20;
	qsin_lut[2458] =  9'sd95;
	icos_lut[2458] = -9'sd39;
	qsin_lut[2459] =  9'sd86;
	icos_lut[2459] = -9'sd57;
	qsin_lut[2460] =  9'sd73;
	icos_lut[2460] = -9'sd73;
	qsin_lut[2461] =  9'sd57;
	icos_lut[2461] = -9'sd86;
	qsin_lut[2462] =  9'sd39;
	icos_lut[2462] = -9'sd95;
	qsin_lut[2463] =  9'sd20;
	icos_lut[2463] = -9'sd101;
	qsin_lut[2464] =  9'sd0;
	icos_lut[2464] = -9'sd101;
	qsin_lut[2465] = -9'sd20;
	icos_lut[2465] = -9'sd99;
	qsin_lut[2466] = -9'sd39;
	icos_lut[2466] = -9'sd93;
	qsin_lut[2467] = -9'sd56;
	icos_lut[2467] = -9'sd84;
	qsin_lut[2468] = -9'sd71;
	icos_lut[2468] = -9'sd71;
	qsin_lut[2469] = -9'sd84;
	icos_lut[2469] = -9'sd56;
	qsin_lut[2470] = -9'sd93;
	icos_lut[2470] = -9'sd39;
	qsin_lut[2471] = -9'sd99;
	icos_lut[2471] = -9'sd20;
	qsin_lut[2472] = -9'sd101;
	icos_lut[2472] = -9'sd0;
	qsin_lut[2473] = -9'sd99;
	icos_lut[2473] =  9'sd20;
	qsin_lut[2474] = -9'sd93;
	icos_lut[2474] =  9'sd39;
	qsin_lut[2475] = -9'sd84;
	icos_lut[2475] =  9'sd56;
	qsin_lut[2476] = -9'sd71;
	icos_lut[2476] =  9'sd71;
	qsin_lut[2477] = -9'sd56;
	icos_lut[2477] =  9'sd84;
	qsin_lut[2478] = -9'sd39;
	icos_lut[2478] =  9'sd93;
	qsin_lut[2479] = -9'sd20;
	icos_lut[2479] =  9'sd99;
	qsin_lut[2480] = -9'sd0;
	icos_lut[2480] =  9'sd101;
	qsin_lut[2481] =  9'sd20;
	icos_lut[2481] =  9'sd99;
	qsin_lut[2482] =  9'sd39;
	icos_lut[2482] =  9'sd93;
	qsin_lut[2483] =  9'sd56;
	icos_lut[2483] =  9'sd84;
	qsin_lut[2484] =  9'sd71;
	icos_lut[2484] =  9'sd71;
	qsin_lut[2485] =  9'sd84;
	icos_lut[2485] =  9'sd56;
	qsin_lut[2486] =  9'sd93;
	icos_lut[2486] =  9'sd39;
	qsin_lut[2487] =  9'sd99;
	icos_lut[2487] =  9'sd20;
	qsin_lut[2488] =  9'sd101;
	icos_lut[2488] =  9'sd0;
	qsin_lut[2489] =  9'sd99;
	icos_lut[2489] = -9'sd20;
	qsin_lut[2490] =  9'sd93;
	icos_lut[2490] = -9'sd39;
	qsin_lut[2491] =  9'sd84;
	icos_lut[2491] = -9'sd56;
	qsin_lut[2492] =  9'sd71;
	icos_lut[2492] = -9'sd71;
	qsin_lut[2493] =  9'sd56;
	icos_lut[2493] = -9'sd84;
	qsin_lut[2494] =  9'sd39;
	icos_lut[2494] = -9'sd93;
	qsin_lut[2495] =  9'sd20;
	icos_lut[2495] = -9'sd99;
	qsin_lut[2496] =  9'sd0;
	icos_lut[2496] = -9'sd99;
	qsin_lut[2497] = -9'sd19;
	icos_lut[2497] = -9'sd97;
	qsin_lut[2498] = -9'sd38;
	icos_lut[2498] = -9'sd91;
	qsin_lut[2499] = -9'sd55;
	icos_lut[2499] = -9'sd82;
	qsin_lut[2500] = -9'sd70;
	icos_lut[2500] = -9'sd70;
	qsin_lut[2501] = -9'sd82;
	icos_lut[2501] = -9'sd55;
	qsin_lut[2502] = -9'sd91;
	icos_lut[2502] = -9'sd38;
	qsin_lut[2503] = -9'sd97;
	icos_lut[2503] = -9'sd19;
	qsin_lut[2504] = -9'sd99;
	icos_lut[2504] = -9'sd0;
	qsin_lut[2505] = -9'sd97;
	icos_lut[2505] =  9'sd19;
	qsin_lut[2506] = -9'sd91;
	icos_lut[2506] =  9'sd38;
	qsin_lut[2507] = -9'sd82;
	icos_lut[2507] =  9'sd55;
	qsin_lut[2508] = -9'sd70;
	icos_lut[2508] =  9'sd70;
	qsin_lut[2509] = -9'sd55;
	icos_lut[2509] =  9'sd82;
	qsin_lut[2510] = -9'sd38;
	icos_lut[2510] =  9'sd91;
	qsin_lut[2511] = -9'sd19;
	icos_lut[2511] =  9'sd97;
	qsin_lut[2512] = -9'sd0;
	icos_lut[2512] =  9'sd99;
	qsin_lut[2513] =  9'sd19;
	icos_lut[2513] =  9'sd97;
	qsin_lut[2514] =  9'sd38;
	icos_lut[2514] =  9'sd91;
	qsin_lut[2515] =  9'sd55;
	icos_lut[2515] =  9'sd82;
	qsin_lut[2516] =  9'sd70;
	icos_lut[2516] =  9'sd70;
	qsin_lut[2517] =  9'sd82;
	icos_lut[2517] =  9'sd55;
	qsin_lut[2518] =  9'sd91;
	icos_lut[2518] =  9'sd38;
	qsin_lut[2519] =  9'sd97;
	icos_lut[2519] =  9'sd19;
	qsin_lut[2520] =  9'sd99;
	icos_lut[2520] =  9'sd0;
	qsin_lut[2521] =  9'sd97;
	icos_lut[2521] = -9'sd19;
	qsin_lut[2522] =  9'sd91;
	icos_lut[2522] = -9'sd38;
	qsin_lut[2523] =  9'sd82;
	icos_lut[2523] = -9'sd55;
	qsin_lut[2524] =  9'sd70;
	icos_lut[2524] = -9'sd70;
	qsin_lut[2525] =  9'sd55;
	icos_lut[2525] = -9'sd82;
	qsin_lut[2526] =  9'sd38;
	icos_lut[2526] = -9'sd91;
	qsin_lut[2527] =  9'sd19;
	icos_lut[2527] = -9'sd97;
	qsin_lut[2528] =  9'sd0;
	icos_lut[2528] = -9'sd97;
	qsin_lut[2529] = -9'sd19;
	icos_lut[2529] = -9'sd95;
	qsin_lut[2530] = -9'sd37;
	icos_lut[2530] = -9'sd90;
	qsin_lut[2531] = -9'sd54;
	icos_lut[2531] = -9'sd81;
	qsin_lut[2532] = -9'sd69;
	icos_lut[2532] = -9'sd69;
	qsin_lut[2533] = -9'sd81;
	icos_lut[2533] = -9'sd54;
	qsin_lut[2534] = -9'sd90;
	icos_lut[2534] = -9'sd37;
	qsin_lut[2535] = -9'sd95;
	icos_lut[2535] = -9'sd19;
	qsin_lut[2536] = -9'sd97;
	icos_lut[2536] = -9'sd0;
	qsin_lut[2537] = -9'sd95;
	icos_lut[2537] =  9'sd19;
	qsin_lut[2538] = -9'sd90;
	icos_lut[2538] =  9'sd37;
	qsin_lut[2539] = -9'sd81;
	icos_lut[2539] =  9'sd54;
	qsin_lut[2540] = -9'sd69;
	icos_lut[2540] =  9'sd69;
	qsin_lut[2541] = -9'sd54;
	icos_lut[2541] =  9'sd81;
	qsin_lut[2542] = -9'sd37;
	icos_lut[2542] =  9'sd90;
	qsin_lut[2543] = -9'sd19;
	icos_lut[2543] =  9'sd95;
	qsin_lut[2544] = -9'sd0;
	icos_lut[2544] =  9'sd97;
	qsin_lut[2545] =  9'sd19;
	icos_lut[2545] =  9'sd95;
	qsin_lut[2546] =  9'sd37;
	icos_lut[2546] =  9'sd90;
	qsin_lut[2547] =  9'sd54;
	icos_lut[2547] =  9'sd81;
	qsin_lut[2548] =  9'sd69;
	icos_lut[2548] =  9'sd69;
	qsin_lut[2549] =  9'sd81;
	icos_lut[2549] =  9'sd54;
	qsin_lut[2550] =  9'sd90;
	icos_lut[2550] =  9'sd37;
	qsin_lut[2551] =  9'sd95;
	icos_lut[2551] =  9'sd19;
	qsin_lut[2552] =  9'sd97;
	icos_lut[2552] =  9'sd0;
	qsin_lut[2553] =  9'sd95;
	icos_lut[2553] = -9'sd19;
	qsin_lut[2554] =  9'sd90;
	icos_lut[2554] = -9'sd37;
	qsin_lut[2555] =  9'sd81;
	icos_lut[2555] = -9'sd54;
	qsin_lut[2556] =  9'sd69;
	icos_lut[2556] = -9'sd69;
	qsin_lut[2557] =  9'sd54;
	icos_lut[2557] = -9'sd81;
	qsin_lut[2558] =  9'sd37;
	icos_lut[2558] = -9'sd90;
	qsin_lut[2559] =  9'sd19;
	icos_lut[2559] = -9'sd95;
	qsin_lut[2560] =  9'sd0;
	icos_lut[2560] = -9'sd95;
	qsin_lut[2561] = -9'sd19;
	icos_lut[2561] = -9'sd93;
	qsin_lut[2562] = -9'sd36;
	icos_lut[2562] = -9'sd88;
	qsin_lut[2563] = -9'sd53;
	icos_lut[2563] = -9'sd79;
	qsin_lut[2564] = -9'sd67;
	icos_lut[2564] = -9'sd67;
	qsin_lut[2565] = -9'sd79;
	icos_lut[2565] = -9'sd53;
	qsin_lut[2566] = -9'sd88;
	icos_lut[2566] = -9'sd36;
	qsin_lut[2567] = -9'sd93;
	icos_lut[2567] = -9'sd19;
	qsin_lut[2568] = -9'sd95;
	icos_lut[2568] = -9'sd0;
	qsin_lut[2569] = -9'sd93;
	icos_lut[2569] =  9'sd19;
	qsin_lut[2570] = -9'sd88;
	icos_lut[2570] =  9'sd36;
	qsin_lut[2571] = -9'sd79;
	icos_lut[2571] =  9'sd53;
	qsin_lut[2572] = -9'sd67;
	icos_lut[2572] =  9'sd67;
	qsin_lut[2573] = -9'sd53;
	icos_lut[2573] =  9'sd79;
	qsin_lut[2574] = -9'sd36;
	icos_lut[2574] =  9'sd88;
	qsin_lut[2575] = -9'sd19;
	icos_lut[2575] =  9'sd93;
	qsin_lut[2576] = -9'sd0;
	icos_lut[2576] =  9'sd95;
	qsin_lut[2577] =  9'sd19;
	icos_lut[2577] =  9'sd93;
	qsin_lut[2578] =  9'sd36;
	icos_lut[2578] =  9'sd88;
	qsin_lut[2579] =  9'sd53;
	icos_lut[2579] =  9'sd79;
	qsin_lut[2580] =  9'sd67;
	icos_lut[2580] =  9'sd67;
	qsin_lut[2581] =  9'sd79;
	icos_lut[2581] =  9'sd53;
	qsin_lut[2582] =  9'sd88;
	icos_lut[2582] =  9'sd36;
	qsin_lut[2583] =  9'sd93;
	icos_lut[2583] =  9'sd19;
	qsin_lut[2584] =  9'sd95;
	icos_lut[2584] =  9'sd0;
	qsin_lut[2585] =  9'sd93;
	icos_lut[2585] = -9'sd19;
	qsin_lut[2586] =  9'sd88;
	icos_lut[2586] = -9'sd36;
	qsin_lut[2587] =  9'sd79;
	icos_lut[2587] = -9'sd53;
	qsin_lut[2588] =  9'sd67;
	icos_lut[2588] = -9'sd67;
	qsin_lut[2589] =  9'sd53;
	icos_lut[2589] = -9'sd79;
	qsin_lut[2590] =  9'sd36;
	icos_lut[2590] = -9'sd88;
	qsin_lut[2591] =  9'sd19;
	icos_lut[2591] = -9'sd93;
	qsin_lut[2592] =  9'sd0;
	icos_lut[2592] = -9'sd93;
	qsin_lut[2593] = -9'sd18;
	icos_lut[2593] = -9'sd91;
	qsin_lut[2594] = -9'sd36;
	icos_lut[2594] = -9'sd86;
	qsin_lut[2595] = -9'sd52;
	icos_lut[2595] = -9'sd77;
	qsin_lut[2596] = -9'sd66;
	icos_lut[2596] = -9'sd66;
	qsin_lut[2597] = -9'sd77;
	icos_lut[2597] = -9'sd52;
	qsin_lut[2598] = -9'sd86;
	icos_lut[2598] = -9'sd36;
	qsin_lut[2599] = -9'sd91;
	icos_lut[2599] = -9'sd18;
	qsin_lut[2600] = -9'sd93;
	icos_lut[2600] = -9'sd0;
	qsin_lut[2601] = -9'sd91;
	icos_lut[2601] =  9'sd18;
	qsin_lut[2602] = -9'sd86;
	icos_lut[2602] =  9'sd36;
	qsin_lut[2603] = -9'sd77;
	icos_lut[2603] =  9'sd52;
	qsin_lut[2604] = -9'sd66;
	icos_lut[2604] =  9'sd66;
	qsin_lut[2605] = -9'sd52;
	icos_lut[2605] =  9'sd77;
	qsin_lut[2606] = -9'sd36;
	icos_lut[2606] =  9'sd86;
	qsin_lut[2607] = -9'sd18;
	icos_lut[2607] =  9'sd91;
	qsin_lut[2608] = -9'sd0;
	icos_lut[2608] =  9'sd93;
	qsin_lut[2609] =  9'sd18;
	icos_lut[2609] =  9'sd91;
	qsin_lut[2610] =  9'sd36;
	icos_lut[2610] =  9'sd86;
	qsin_lut[2611] =  9'sd52;
	icos_lut[2611] =  9'sd77;
	qsin_lut[2612] =  9'sd66;
	icos_lut[2612] =  9'sd66;
	qsin_lut[2613] =  9'sd77;
	icos_lut[2613] =  9'sd52;
	qsin_lut[2614] =  9'sd86;
	icos_lut[2614] =  9'sd36;
	qsin_lut[2615] =  9'sd91;
	icos_lut[2615] =  9'sd18;
	qsin_lut[2616] =  9'sd93;
	icos_lut[2616] =  9'sd0;
	qsin_lut[2617] =  9'sd91;
	icos_lut[2617] = -9'sd18;
	qsin_lut[2618] =  9'sd86;
	icos_lut[2618] = -9'sd36;
	qsin_lut[2619] =  9'sd77;
	icos_lut[2619] = -9'sd52;
	qsin_lut[2620] =  9'sd66;
	icos_lut[2620] = -9'sd66;
	qsin_lut[2621] =  9'sd52;
	icos_lut[2621] = -9'sd77;
	qsin_lut[2622] =  9'sd36;
	icos_lut[2622] = -9'sd86;
	qsin_lut[2623] =  9'sd18;
	icos_lut[2623] = -9'sd91;
	qsin_lut[2624] =  9'sd0;
	icos_lut[2624] = -9'sd91;
	qsin_lut[2625] = -9'sd18;
	icos_lut[2625] = -9'sd89;
	qsin_lut[2626] = -9'sd35;
	icos_lut[2626] = -9'sd84;
	qsin_lut[2627] = -9'sd51;
	icos_lut[2627] = -9'sd76;
	qsin_lut[2628] = -9'sd64;
	icos_lut[2628] = -9'sd64;
	qsin_lut[2629] = -9'sd76;
	icos_lut[2629] = -9'sd51;
	qsin_lut[2630] = -9'sd84;
	icos_lut[2630] = -9'sd35;
	qsin_lut[2631] = -9'sd89;
	icos_lut[2631] = -9'sd18;
	qsin_lut[2632] = -9'sd91;
	icos_lut[2632] = -9'sd0;
	qsin_lut[2633] = -9'sd89;
	icos_lut[2633] =  9'sd18;
	qsin_lut[2634] = -9'sd84;
	icos_lut[2634] =  9'sd35;
	qsin_lut[2635] = -9'sd76;
	icos_lut[2635] =  9'sd51;
	qsin_lut[2636] = -9'sd64;
	icos_lut[2636] =  9'sd64;
	qsin_lut[2637] = -9'sd51;
	icos_lut[2637] =  9'sd76;
	qsin_lut[2638] = -9'sd35;
	icos_lut[2638] =  9'sd84;
	qsin_lut[2639] = -9'sd18;
	icos_lut[2639] =  9'sd89;
	qsin_lut[2640] = -9'sd0;
	icos_lut[2640] =  9'sd91;
	qsin_lut[2641] =  9'sd18;
	icos_lut[2641] =  9'sd89;
	qsin_lut[2642] =  9'sd35;
	icos_lut[2642] =  9'sd84;
	qsin_lut[2643] =  9'sd51;
	icos_lut[2643] =  9'sd76;
	qsin_lut[2644] =  9'sd64;
	icos_lut[2644] =  9'sd64;
	qsin_lut[2645] =  9'sd76;
	icos_lut[2645] =  9'sd51;
	qsin_lut[2646] =  9'sd84;
	icos_lut[2646] =  9'sd35;
	qsin_lut[2647] =  9'sd89;
	icos_lut[2647] =  9'sd18;
	qsin_lut[2648] =  9'sd91;
	icos_lut[2648] =  9'sd0;
	qsin_lut[2649] =  9'sd89;
	icos_lut[2649] = -9'sd18;
	qsin_lut[2650] =  9'sd84;
	icos_lut[2650] = -9'sd35;
	qsin_lut[2651] =  9'sd76;
	icos_lut[2651] = -9'sd51;
	qsin_lut[2652] =  9'sd64;
	icos_lut[2652] = -9'sd64;
	qsin_lut[2653] =  9'sd51;
	icos_lut[2653] = -9'sd76;
	qsin_lut[2654] =  9'sd35;
	icos_lut[2654] = -9'sd84;
	qsin_lut[2655] =  9'sd18;
	icos_lut[2655] = -9'sd89;
	qsin_lut[2656] =  9'sd0;
	icos_lut[2656] = -9'sd89;
	qsin_lut[2657] = -9'sd17;
	icos_lut[2657] = -9'sd87;
	qsin_lut[2658] = -9'sd34;
	icos_lut[2658] = -9'sd82;
	qsin_lut[2659] = -9'sd49;
	icos_lut[2659] = -9'sd74;
	qsin_lut[2660] = -9'sd63;
	icos_lut[2660] = -9'sd63;
	qsin_lut[2661] = -9'sd74;
	icos_lut[2661] = -9'sd49;
	qsin_lut[2662] = -9'sd82;
	icos_lut[2662] = -9'sd34;
	qsin_lut[2663] = -9'sd87;
	icos_lut[2663] = -9'sd17;
	qsin_lut[2664] = -9'sd89;
	icos_lut[2664] = -9'sd0;
	qsin_lut[2665] = -9'sd87;
	icos_lut[2665] =  9'sd17;
	qsin_lut[2666] = -9'sd82;
	icos_lut[2666] =  9'sd34;
	qsin_lut[2667] = -9'sd74;
	icos_lut[2667] =  9'sd49;
	qsin_lut[2668] = -9'sd63;
	icos_lut[2668] =  9'sd63;
	qsin_lut[2669] = -9'sd49;
	icos_lut[2669] =  9'sd74;
	qsin_lut[2670] = -9'sd34;
	icos_lut[2670] =  9'sd82;
	qsin_lut[2671] = -9'sd17;
	icos_lut[2671] =  9'sd87;
	qsin_lut[2672] = -9'sd0;
	icos_lut[2672] =  9'sd89;
	qsin_lut[2673] =  9'sd17;
	icos_lut[2673] =  9'sd87;
	qsin_lut[2674] =  9'sd34;
	icos_lut[2674] =  9'sd82;
	qsin_lut[2675] =  9'sd49;
	icos_lut[2675] =  9'sd74;
	qsin_lut[2676] =  9'sd63;
	icos_lut[2676] =  9'sd63;
	qsin_lut[2677] =  9'sd74;
	icos_lut[2677] =  9'sd49;
	qsin_lut[2678] =  9'sd82;
	icos_lut[2678] =  9'sd34;
	qsin_lut[2679] =  9'sd87;
	icos_lut[2679] =  9'sd17;
	qsin_lut[2680] =  9'sd89;
	icos_lut[2680] =  9'sd0;
	qsin_lut[2681] =  9'sd87;
	icos_lut[2681] = -9'sd17;
	qsin_lut[2682] =  9'sd82;
	icos_lut[2682] = -9'sd34;
	qsin_lut[2683] =  9'sd74;
	icos_lut[2683] = -9'sd49;
	qsin_lut[2684] =  9'sd63;
	icos_lut[2684] = -9'sd63;
	qsin_lut[2685] =  9'sd49;
	icos_lut[2685] = -9'sd74;
	qsin_lut[2686] =  9'sd34;
	icos_lut[2686] = -9'sd82;
	qsin_lut[2687] =  9'sd17;
	icos_lut[2687] = -9'sd87;
	qsin_lut[2688] =  9'sd0;
	icos_lut[2688] = -9'sd87;
	qsin_lut[2689] = -9'sd17;
	icos_lut[2689] = -9'sd85;
	qsin_lut[2690] = -9'sd33;
	icos_lut[2690] = -9'sd80;
	qsin_lut[2691] = -9'sd48;
	icos_lut[2691] = -9'sd72;
	qsin_lut[2692] = -9'sd62;
	icos_lut[2692] = -9'sd62;
	qsin_lut[2693] = -9'sd72;
	icos_lut[2693] = -9'sd48;
	qsin_lut[2694] = -9'sd80;
	icos_lut[2694] = -9'sd33;
	qsin_lut[2695] = -9'sd85;
	icos_lut[2695] = -9'sd17;
	qsin_lut[2696] = -9'sd87;
	icos_lut[2696] = -9'sd0;
	qsin_lut[2697] = -9'sd85;
	icos_lut[2697] =  9'sd17;
	qsin_lut[2698] = -9'sd80;
	icos_lut[2698] =  9'sd33;
	qsin_lut[2699] = -9'sd72;
	icos_lut[2699] =  9'sd48;
	qsin_lut[2700] = -9'sd62;
	icos_lut[2700] =  9'sd62;
	qsin_lut[2701] = -9'sd48;
	icos_lut[2701] =  9'sd72;
	qsin_lut[2702] = -9'sd33;
	icos_lut[2702] =  9'sd80;
	qsin_lut[2703] = -9'sd17;
	icos_lut[2703] =  9'sd85;
	qsin_lut[2704] = -9'sd0;
	icos_lut[2704] =  9'sd87;
	qsin_lut[2705] =  9'sd17;
	icos_lut[2705] =  9'sd85;
	qsin_lut[2706] =  9'sd33;
	icos_lut[2706] =  9'sd80;
	qsin_lut[2707] =  9'sd48;
	icos_lut[2707] =  9'sd72;
	qsin_lut[2708] =  9'sd62;
	icos_lut[2708] =  9'sd62;
	qsin_lut[2709] =  9'sd72;
	icos_lut[2709] =  9'sd48;
	qsin_lut[2710] =  9'sd80;
	icos_lut[2710] =  9'sd33;
	qsin_lut[2711] =  9'sd85;
	icos_lut[2711] =  9'sd17;
	qsin_lut[2712] =  9'sd87;
	icos_lut[2712] =  9'sd0;
	qsin_lut[2713] =  9'sd85;
	icos_lut[2713] = -9'sd17;
	qsin_lut[2714] =  9'sd80;
	icos_lut[2714] = -9'sd33;
	qsin_lut[2715] =  9'sd72;
	icos_lut[2715] = -9'sd48;
	qsin_lut[2716] =  9'sd62;
	icos_lut[2716] = -9'sd62;
	qsin_lut[2717] =  9'sd48;
	icos_lut[2717] = -9'sd72;
	qsin_lut[2718] =  9'sd33;
	icos_lut[2718] = -9'sd80;
	qsin_lut[2719] =  9'sd17;
	icos_lut[2719] = -9'sd85;
	qsin_lut[2720] =  9'sd0;
	icos_lut[2720] = -9'sd85;
	qsin_lut[2721] = -9'sd17;
	icos_lut[2721] = -9'sd83;
	qsin_lut[2722] = -9'sd33;
	icos_lut[2722] = -9'sd79;
	qsin_lut[2723] = -9'sd47;
	icos_lut[2723] = -9'sd71;
	qsin_lut[2724] = -9'sd60;
	icos_lut[2724] = -9'sd60;
	qsin_lut[2725] = -9'sd71;
	icos_lut[2725] = -9'sd47;
	qsin_lut[2726] = -9'sd79;
	icos_lut[2726] = -9'sd33;
	qsin_lut[2727] = -9'sd83;
	icos_lut[2727] = -9'sd17;
	qsin_lut[2728] = -9'sd85;
	icos_lut[2728] = -9'sd0;
	qsin_lut[2729] = -9'sd83;
	icos_lut[2729] =  9'sd17;
	qsin_lut[2730] = -9'sd79;
	icos_lut[2730] =  9'sd33;
	qsin_lut[2731] = -9'sd71;
	icos_lut[2731] =  9'sd47;
	qsin_lut[2732] = -9'sd60;
	icos_lut[2732] =  9'sd60;
	qsin_lut[2733] = -9'sd47;
	icos_lut[2733] =  9'sd71;
	qsin_lut[2734] = -9'sd33;
	icos_lut[2734] =  9'sd79;
	qsin_lut[2735] = -9'sd17;
	icos_lut[2735] =  9'sd83;
	qsin_lut[2736] = -9'sd0;
	icos_lut[2736] =  9'sd85;
	qsin_lut[2737] =  9'sd17;
	icos_lut[2737] =  9'sd83;
	qsin_lut[2738] =  9'sd33;
	icos_lut[2738] =  9'sd79;
	qsin_lut[2739] =  9'sd47;
	icos_lut[2739] =  9'sd71;
	qsin_lut[2740] =  9'sd60;
	icos_lut[2740] =  9'sd60;
	qsin_lut[2741] =  9'sd71;
	icos_lut[2741] =  9'sd47;
	qsin_lut[2742] =  9'sd79;
	icos_lut[2742] =  9'sd33;
	qsin_lut[2743] =  9'sd83;
	icos_lut[2743] =  9'sd17;
	qsin_lut[2744] =  9'sd85;
	icos_lut[2744] =  9'sd0;
	qsin_lut[2745] =  9'sd83;
	icos_lut[2745] = -9'sd17;
	qsin_lut[2746] =  9'sd79;
	icos_lut[2746] = -9'sd33;
	qsin_lut[2747] =  9'sd71;
	icos_lut[2747] = -9'sd47;
	qsin_lut[2748] =  9'sd60;
	icos_lut[2748] = -9'sd60;
	qsin_lut[2749] =  9'sd47;
	icos_lut[2749] = -9'sd71;
	qsin_lut[2750] =  9'sd33;
	icos_lut[2750] = -9'sd79;
	qsin_lut[2751] =  9'sd17;
	icos_lut[2751] = -9'sd83;
	qsin_lut[2752] =  9'sd0;
	icos_lut[2752] = -9'sd83;
	qsin_lut[2753] = -9'sd16;
	icos_lut[2753] = -9'sd81;
	qsin_lut[2754] = -9'sd32;
	icos_lut[2754] = -9'sd77;
	qsin_lut[2755] = -9'sd46;
	icos_lut[2755] = -9'sd69;
	qsin_lut[2756] = -9'sd59;
	icos_lut[2756] = -9'sd59;
	qsin_lut[2757] = -9'sd69;
	icos_lut[2757] = -9'sd46;
	qsin_lut[2758] = -9'sd77;
	icos_lut[2758] = -9'sd32;
	qsin_lut[2759] = -9'sd81;
	icos_lut[2759] = -9'sd16;
	qsin_lut[2760] = -9'sd83;
	icos_lut[2760] = -9'sd0;
	qsin_lut[2761] = -9'sd81;
	icos_lut[2761] =  9'sd16;
	qsin_lut[2762] = -9'sd77;
	icos_lut[2762] =  9'sd32;
	qsin_lut[2763] = -9'sd69;
	icos_lut[2763] =  9'sd46;
	qsin_lut[2764] = -9'sd59;
	icos_lut[2764] =  9'sd59;
	qsin_lut[2765] = -9'sd46;
	icos_lut[2765] =  9'sd69;
	qsin_lut[2766] = -9'sd32;
	icos_lut[2766] =  9'sd77;
	qsin_lut[2767] = -9'sd16;
	icos_lut[2767] =  9'sd81;
	qsin_lut[2768] = -9'sd0;
	icos_lut[2768] =  9'sd83;
	qsin_lut[2769] =  9'sd16;
	icos_lut[2769] =  9'sd81;
	qsin_lut[2770] =  9'sd32;
	icos_lut[2770] =  9'sd77;
	qsin_lut[2771] =  9'sd46;
	icos_lut[2771] =  9'sd69;
	qsin_lut[2772] =  9'sd59;
	icos_lut[2772] =  9'sd59;
	qsin_lut[2773] =  9'sd69;
	icos_lut[2773] =  9'sd46;
	qsin_lut[2774] =  9'sd77;
	icos_lut[2774] =  9'sd32;
	qsin_lut[2775] =  9'sd81;
	icos_lut[2775] =  9'sd16;
	qsin_lut[2776] =  9'sd83;
	icos_lut[2776] =  9'sd0;
	qsin_lut[2777] =  9'sd81;
	icos_lut[2777] = -9'sd16;
	qsin_lut[2778] =  9'sd77;
	icos_lut[2778] = -9'sd32;
	qsin_lut[2779] =  9'sd69;
	icos_lut[2779] = -9'sd46;
	qsin_lut[2780] =  9'sd59;
	icos_lut[2780] = -9'sd59;
	qsin_lut[2781] =  9'sd46;
	icos_lut[2781] = -9'sd69;
	qsin_lut[2782] =  9'sd32;
	icos_lut[2782] = -9'sd77;
	qsin_lut[2783] =  9'sd16;
	icos_lut[2783] = -9'sd81;
	qsin_lut[2784] =  9'sd0;
	icos_lut[2784] = -9'sd81;
	qsin_lut[2785] = -9'sd16;
	icos_lut[2785] = -9'sd79;
	qsin_lut[2786] = -9'sd31;
	icos_lut[2786] = -9'sd75;
	qsin_lut[2787] = -9'sd45;
	icos_lut[2787] = -9'sd67;
	qsin_lut[2788] = -9'sd57;
	icos_lut[2788] = -9'sd57;
	qsin_lut[2789] = -9'sd67;
	icos_lut[2789] = -9'sd45;
	qsin_lut[2790] = -9'sd75;
	icos_lut[2790] = -9'sd31;
	qsin_lut[2791] = -9'sd79;
	icos_lut[2791] = -9'sd16;
	qsin_lut[2792] = -9'sd81;
	icos_lut[2792] = -9'sd0;
	qsin_lut[2793] = -9'sd79;
	icos_lut[2793] =  9'sd16;
	qsin_lut[2794] = -9'sd75;
	icos_lut[2794] =  9'sd31;
	qsin_lut[2795] = -9'sd67;
	icos_lut[2795] =  9'sd45;
	qsin_lut[2796] = -9'sd57;
	icos_lut[2796] =  9'sd57;
	qsin_lut[2797] = -9'sd45;
	icos_lut[2797] =  9'sd67;
	qsin_lut[2798] = -9'sd31;
	icos_lut[2798] =  9'sd75;
	qsin_lut[2799] = -9'sd16;
	icos_lut[2799] =  9'sd79;
	qsin_lut[2800] = -9'sd0;
	icos_lut[2800] =  9'sd81;
	qsin_lut[2801] =  9'sd16;
	icos_lut[2801] =  9'sd79;
	qsin_lut[2802] =  9'sd31;
	icos_lut[2802] =  9'sd75;
	qsin_lut[2803] =  9'sd45;
	icos_lut[2803] =  9'sd67;
	qsin_lut[2804] =  9'sd57;
	icos_lut[2804] =  9'sd57;
	qsin_lut[2805] =  9'sd67;
	icos_lut[2805] =  9'sd45;
	qsin_lut[2806] =  9'sd75;
	icos_lut[2806] =  9'sd31;
	qsin_lut[2807] =  9'sd79;
	icos_lut[2807] =  9'sd16;
	qsin_lut[2808] =  9'sd81;
	icos_lut[2808] =  9'sd0;
	qsin_lut[2809] =  9'sd79;
	icos_lut[2809] = -9'sd16;
	qsin_lut[2810] =  9'sd75;
	icos_lut[2810] = -9'sd31;
	qsin_lut[2811] =  9'sd67;
	icos_lut[2811] = -9'sd45;
	qsin_lut[2812] =  9'sd57;
	icos_lut[2812] = -9'sd57;
	qsin_lut[2813] =  9'sd45;
	icos_lut[2813] = -9'sd67;
	qsin_lut[2814] =  9'sd31;
	icos_lut[2814] = -9'sd75;
	qsin_lut[2815] =  9'sd16;
	icos_lut[2815] = -9'sd79;
	qsin_lut[2816] =  9'sd0;
	icos_lut[2816] = -9'sd79;
	qsin_lut[2817] = -9'sd15;
	icos_lut[2817] = -9'sd77;
	qsin_lut[2818] = -9'sd30;
	icos_lut[2818] = -9'sd73;
	qsin_lut[2819] = -9'sd44;
	icos_lut[2819] = -9'sd66;
	qsin_lut[2820] = -9'sd56;
	icos_lut[2820] = -9'sd56;
	qsin_lut[2821] = -9'sd66;
	icos_lut[2821] = -9'sd44;
	qsin_lut[2822] = -9'sd73;
	icos_lut[2822] = -9'sd30;
	qsin_lut[2823] = -9'sd77;
	icos_lut[2823] = -9'sd15;
	qsin_lut[2824] = -9'sd79;
	icos_lut[2824] = -9'sd0;
	qsin_lut[2825] = -9'sd77;
	icos_lut[2825] =  9'sd15;
	qsin_lut[2826] = -9'sd73;
	icos_lut[2826] =  9'sd30;
	qsin_lut[2827] = -9'sd66;
	icos_lut[2827] =  9'sd44;
	qsin_lut[2828] = -9'sd56;
	icos_lut[2828] =  9'sd56;
	qsin_lut[2829] = -9'sd44;
	icos_lut[2829] =  9'sd66;
	qsin_lut[2830] = -9'sd30;
	icos_lut[2830] =  9'sd73;
	qsin_lut[2831] = -9'sd15;
	icos_lut[2831] =  9'sd77;
	qsin_lut[2832] = -9'sd0;
	icos_lut[2832] =  9'sd79;
	qsin_lut[2833] =  9'sd15;
	icos_lut[2833] =  9'sd77;
	qsin_lut[2834] =  9'sd30;
	icos_lut[2834] =  9'sd73;
	qsin_lut[2835] =  9'sd44;
	icos_lut[2835] =  9'sd66;
	qsin_lut[2836] =  9'sd56;
	icos_lut[2836] =  9'sd56;
	qsin_lut[2837] =  9'sd66;
	icos_lut[2837] =  9'sd44;
	qsin_lut[2838] =  9'sd73;
	icos_lut[2838] =  9'sd30;
	qsin_lut[2839] =  9'sd77;
	icos_lut[2839] =  9'sd15;
	qsin_lut[2840] =  9'sd79;
	icos_lut[2840] =  9'sd0;
	qsin_lut[2841] =  9'sd77;
	icos_lut[2841] = -9'sd15;
	qsin_lut[2842] =  9'sd73;
	icos_lut[2842] = -9'sd30;
	qsin_lut[2843] =  9'sd66;
	icos_lut[2843] = -9'sd44;
	qsin_lut[2844] =  9'sd56;
	icos_lut[2844] = -9'sd56;
	qsin_lut[2845] =  9'sd44;
	icos_lut[2845] = -9'sd66;
	qsin_lut[2846] =  9'sd30;
	icos_lut[2846] = -9'sd73;
	qsin_lut[2847] =  9'sd15;
	icos_lut[2847] = -9'sd77;
	qsin_lut[2848] =  9'sd0;
	icos_lut[2848] = -9'sd77;
	qsin_lut[2849] = -9'sd15;
	icos_lut[2849] = -9'sd76;
	qsin_lut[2850] = -9'sd29;
	icos_lut[2850] = -9'sd71;
	qsin_lut[2851] = -9'sd43;
	icos_lut[2851] = -9'sd64;
	qsin_lut[2852] = -9'sd54;
	icos_lut[2852] = -9'sd54;
	qsin_lut[2853] = -9'sd64;
	icos_lut[2853] = -9'sd43;
	qsin_lut[2854] = -9'sd71;
	icos_lut[2854] = -9'sd29;
	qsin_lut[2855] = -9'sd76;
	icos_lut[2855] = -9'sd15;
	qsin_lut[2856] = -9'sd77;
	icos_lut[2856] = -9'sd0;
	qsin_lut[2857] = -9'sd76;
	icos_lut[2857] =  9'sd15;
	qsin_lut[2858] = -9'sd71;
	icos_lut[2858] =  9'sd29;
	qsin_lut[2859] = -9'sd64;
	icos_lut[2859] =  9'sd43;
	qsin_lut[2860] = -9'sd54;
	icos_lut[2860] =  9'sd54;
	qsin_lut[2861] = -9'sd43;
	icos_lut[2861] =  9'sd64;
	qsin_lut[2862] = -9'sd29;
	icos_lut[2862] =  9'sd71;
	qsin_lut[2863] = -9'sd15;
	icos_lut[2863] =  9'sd76;
	qsin_lut[2864] = -9'sd0;
	icos_lut[2864] =  9'sd77;
	qsin_lut[2865] =  9'sd15;
	icos_lut[2865] =  9'sd76;
	qsin_lut[2866] =  9'sd29;
	icos_lut[2866] =  9'sd71;
	qsin_lut[2867] =  9'sd43;
	icos_lut[2867] =  9'sd64;
	qsin_lut[2868] =  9'sd54;
	icos_lut[2868] =  9'sd54;
	qsin_lut[2869] =  9'sd64;
	icos_lut[2869] =  9'sd43;
	qsin_lut[2870] =  9'sd71;
	icos_lut[2870] =  9'sd29;
	qsin_lut[2871] =  9'sd76;
	icos_lut[2871] =  9'sd15;
	qsin_lut[2872] =  9'sd77;
	icos_lut[2872] =  9'sd0;
	qsin_lut[2873] =  9'sd76;
	icos_lut[2873] = -9'sd15;
	qsin_lut[2874] =  9'sd71;
	icos_lut[2874] = -9'sd29;
	qsin_lut[2875] =  9'sd64;
	icos_lut[2875] = -9'sd43;
	qsin_lut[2876] =  9'sd54;
	icos_lut[2876] = -9'sd54;
	qsin_lut[2877] =  9'sd43;
	icos_lut[2877] = -9'sd64;
	qsin_lut[2878] =  9'sd29;
	icos_lut[2878] = -9'sd71;
	qsin_lut[2879] =  9'sd15;
	icos_lut[2879] = -9'sd76;
	qsin_lut[2880] =  9'sd0;
	icos_lut[2880] = -9'sd75;
	qsin_lut[2881] = -9'sd15;
	icos_lut[2881] = -9'sd74;
	qsin_lut[2882] = -9'sd29;
	icos_lut[2882] = -9'sd69;
	qsin_lut[2883] = -9'sd42;
	icos_lut[2883] = -9'sd62;
	qsin_lut[2884] = -9'sd53;
	icos_lut[2884] = -9'sd53;
	qsin_lut[2885] = -9'sd62;
	icos_lut[2885] = -9'sd42;
	qsin_lut[2886] = -9'sd69;
	icos_lut[2886] = -9'sd29;
	qsin_lut[2887] = -9'sd74;
	icos_lut[2887] = -9'sd15;
	qsin_lut[2888] = -9'sd75;
	icos_lut[2888] = -9'sd0;
	qsin_lut[2889] = -9'sd74;
	icos_lut[2889] =  9'sd15;
	qsin_lut[2890] = -9'sd69;
	icos_lut[2890] =  9'sd29;
	qsin_lut[2891] = -9'sd62;
	icos_lut[2891] =  9'sd42;
	qsin_lut[2892] = -9'sd53;
	icos_lut[2892] =  9'sd53;
	qsin_lut[2893] = -9'sd42;
	icos_lut[2893] =  9'sd62;
	qsin_lut[2894] = -9'sd29;
	icos_lut[2894] =  9'sd69;
	qsin_lut[2895] = -9'sd15;
	icos_lut[2895] =  9'sd74;
	qsin_lut[2896] = -9'sd0;
	icos_lut[2896] =  9'sd75;
	qsin_lut[2897] =  9'sd15;
	icos_lut[2897] =  9'sd74;
	qsin_lut[2898] =  9'sd29;
	icos_lut[2898] =  9'sd69;
	qsin_lut[2899] =  9'sd42;
	icos_lut[2899] =  9'sd62;
	qsin_lut[2900] =  9'sd53;
	icos_lut[2900] =  9'sd53;
	qsin_lut[2901] =  9'sd62;
	icos_lut[2901] =  9'sd42;
	qsin_lut[2902] =  9'sd69;
	icos_lut[2902] =  9'sd29;
	qsin_lut[2903] =  9'sd74;
	icos_lut[2903] =  9'sd15;
	qsin_lut[2904] =  9'sd75;
	icos_lut[2904] =  9'sd0;
	qsin_lut[2905] =  9'sd74;
	icos_lut[2905] = -9'sd15;
	qsin_lut[2906] =  9'sd69;
	icos_lut[2906] = -9'sd29;
	qsin_lut[2907] =  9'sd62;
	icos_lut[2907] = -9'sd42;
	qsin_lut[2908] =  9'sd53;
	icos_lut[2908] = -9'sd53;
	qsin_lut[2909] =  9'sd42;
	icos_lut[2909] = -9'sd62;
	qsin_lut[2910] =  9'sd29;
	icos_lut[2910] = -9'sd69;
	qsin_lut[2911] =  9'sd15;
	icos_lut[2911] = -9'sd74;
	qsin_lut[2912] =  9'sd0;
	icos_lut[2912] = -9'sd73;
	qsin_lut[2913] = -9'sd14;
	icos_lut[2913] = -9'sd72;
	qsin_lut[2914] = -9'sd28;
	icos_lut[2914] = -9'sd67;
	qsin_lut[2915] = -9'sd41;
	icos_lut[2915] = -9'sd61;
	qsin_lut[2916] = -9'sd52;
	icos_lut[2916] = -9'sd52;
	qsin_lut[2917] = -9'sd61;
	icos_lut[2917] = -9'sd41;
	qsin_lut[2918] = -9'sd67;
	icos_lut[2918] = -9'sd28;
	qsin_lut[2919] = -9'sd72;
	icos_lut[2919] = -9'sd14;
	qsin_lut[2920] = -9'sd73;
	icos_lut[2920] = -9'sd0;
	qsin_lut[2921] = -9'sd72;
	icos_lut[2921] =  9'sd14;
	qsin_lut[2922] = -9'sd67;
	icos_lut[2922] =  9'sd28;
	qsin_lut[2923] = -9'sd61;
	icos_lut[2923] =  9'sd41;
	qsin_lut[2924] = -9'sd52;
	icos_lut[2924] =  9'sd52;
	qsin_lut[2925] = -9'sd41;
	icos_lut[2925] =  9'sd61;
	qsin_lut[2926] = -9'sd28;
	icos_lut[2926] =  9'sd67;
	qsin_lut[2927] = -9'sd14;
	icos_lut[2927] =  9'sd72;
	qsin_lut[2928] = -9'sd0;
	icos_lut[2928] =  9'sd73;
	qsin_lut[2929] =  9'sd14;
	icos_lut[2929] =  9'sd72;
	qsin_lut[2930] =  9'sd28;
	icos_lut[2930] =  9'sd67;
	qsin_lut[2931] =  9'sd41;
	icos_lut[2931] =  9'sd61;
	qsin_lut[2932] =  9'sd52;
	icos_lut[2932] =  9'sd52;
	qsin_lut[2933] =  9'sd61;
	icos_lut[2933] =  9'sd41;
	qsin_lut[2934] =  9'sd67;
	icos_lut[2934] =  9'sd28;
	qsin_lut[2935] =  9'sd72;
	icos_lut[2935] =  9'sd14;
	qsin_lut[2936] =  9'sd73;
	icos_lut[2936] =  9'sd0;
	qsin_lut[2937] =  9'sd72;
	icos_lut[2937] = -9'sd14;
	qsin_lut[2938] =  9'sd67;
	icos_lut[2938] = -9'sd28;
	qsin_lut[2939] =  9'sd61;
	icos_lut[2939] = -9'sd41;
	qsin_lut[2940] =  9'sd52;
	icos_lut[2940] = -9'sd52;
	qsin_lut[2941] =  9'sd41;
	icos_lut[2941] = -9'sd61;
	qsin_lut[2942] =  9'sd28;
	icos_lut[2942] = -9'sd67;
	qsin_lut[2943] =  9'sd14;
	icos_lut[2943] = -9'sd72;
	qsin_lut[2944] =  9'sd0;
	icos_lut[2944] = -9'sd71;
	qsin_lut[2945] = -9'sd14;
	icos_lut[2945] = -9'sd70;
	qsin_lut[2946] = -9'sd27;
	icos_lut[2946] = -9'sd66;
	qsin_lut[2947] = -9'sd39;
	icos_lut[2947] = -9'sd59;
	qsin_lut[2948] = -9'sd50;
	icos_lut[2948] = -9'sd50;
	qsin_lut[2949] = -9'sd59;
	icos_lut[2949] = -9'sd39;
	qsin_lut[2950] = -9'sd66;
	icos_lut[2950] = -9'sd27;
	qsin_lut[2951] = -9'sd70;
	icos_lut[2951] = -9'sd14;
	qsin_lut[2952] = -9'sd71;
	icos_lut[2952] = -9'sd0;
	qsin_lut[2953] = -9'sd70;
	icos_lut[2953] =  9'sd14;
	qsin_lut[2954] = -9'sd66;
	icos_lut[2954] =  9'sd27;
	qsin_lut[2955] = -9'sd59;
	icos_lut[2955] =  9'sd39;
	qsin_lut[2956] = -9'sd50;
	icos_lut[2956] =  9'sd50;
	qsin_lut[2957] = -9'sd39;
	icos_lut[2957] =  9'sd59;
	qsin_lut[2958] = -9'sd27;
	icos_lut[2958] =  9'sd66;
	qsin_lut[2959] = -9'sd14;
	icos_lut[2959] =  9'sd70;
	qsin_lut[2960] = -9'sd0;
	icos_lut[2960] =  9'sd71;
	qsin_lut[2961] =  9'sd14;
	icos_lut[2961] =  9'sd70;
	qsin_lut[2962] =  9'sd27;
	icos_lut[2962] =  9'sd66;
	qsin_lut[2963] =  9'sd39;
	icos_lut[2963] =  9'sd59;
	qsin_lut[2964] =  9'sd50;
	icos_lut[2964] =  9'sd50;
	qsin_lut[2965] =  9'sd59;
	icos_lut[2965] =  9'sd39;
	qsin_lut[2966] =  9'sd66;
	icos_lut[2966] =  9'sd27;
	qsin_lut[2967] =  9'sd70;
	icos_lut[2967] =  9'sd14;
	qsin_lut[2968] =  9'sd71;
	icos_lut[2968] =  9'sd0;
	qsin_lut[2969] =  9'sd70;
	icos_lut[2969] = -9'sd14;
	qsin_lut[2970] =  9'sd66;
	icos_lut[2970] = -9'sd27;
	qsin_lut[2971] =  9'sd59;
	icos_lut[2971] = -9'sd39;
	qsin_lut[2972] =  9'sd50;
	icos_lut[2972] = -9'sd50;
	qsin_lut[2973] =  9'sd39;
	icos_lut[2973] = -9'sd59;
	qsin_lut[2974] =  9'sd27;
	icos_lut[2974] = -9'sd66;
	qsin_lut[2975] =  9'sd14;
	icos_lut[2975] = -9'sd70;
	qsin_lut[2976] =  9'sd0;
	icos_lut[2976] = -9'sd69;
	qsin_lut[2977] = -9'sd13;
	icos_lut[2977] = -9'sd68;
	qsin_lut[2978] = -9'sd26;
	icos_lut[2978] = -9'sd64;
	qsin_lut[2979] = -9'sd38;
	icos_lut[2979] = -9'sd57;
	qsin_lut[2980] = -9'sd49;
	icos_lut[2980] = -9'sd49;
	qsin_lut[2981] = -9'sd57;
	icos_lut[2981] = -9'sd38;
	qsin_lut[2982] = -9'sd64;
	icos_lut[2982] = -9'sd26;
	qsin_lut[2983] = -9'sd68;
	icos_lut[2983] = -9'sd13;
	qsin_lut[2984] = -9'sd69;
	icos_lut[2984] = -9'sd0;
	qsin_lut[2985] = -9'sd68;
	icos_lut[2985] =  9'sd13;
	qsin_lut[2986] = -9'sd64;
	icos_lut[2986] =  9'sd26;
	qsin_lut[2987] = -9'sd57;
	icos_lut[2987] =  9'sd38;
	qsin_lut[2988] = -9'sd49;
	icos_lut[2988] =  9'sd49;
	qsin_lut[2989] = -9'sd38;
	icos_lut[2989] =  9'sd57;
	qsin_lut[2990] = -9'sd26;
	icos_lut[2990] =  9'sd64;
	qsin_lut[2991] = -9'sd13;
	icos_lut[2991] =  9'sd68;
	qsin_lut[2992] = -9'sd0;
	icos_lut[2992] =  9'sd69;
	qsin_lut[2993] =  9'sd13;
	icos_lut[2993] =  9'sd68;
	qsin_lut[2994] =  9'sd26;
	icos_lut[2994] =  9'sd64;
	qsin_lut[2995] =  9'sd38;
	icos_lut[2995] =  9'sd57;
	qsin_lut[2996] =  9'sd49;
	icos_lut[2996] =  9'sd49;
	qsin_lut[2997] =  9'sd57;
	icos_lut[2997] =  9'sd38;
	qsin_lut[2998] =  9'sd64;
	icos_lut[2998] =  9'sd26;
	qsin_lut[2999] =  9'sd68;
	icos_lut[2999] =  9'sd13;
	qsin_lut[3000] =  9'sd69;
	icos_lut[3000] =  9'sd0;
	qsin_lut[3001] =  9'sd68;
	icos_lut[3001] = -9'sd13;
	qsin_lut[3002] =  9'sd64;
	icos_lut[3002] = -9'sd26;
	qsin_lut[3003] =  9'sd57;
	icos_lut[3003] = -9'sd38;
	qsin_lut[3004] =  9'sd49;
	icos_lut[3004] = -9'sd49;
	qsin_lut[3005] =  9'sd38;
	icos_lut[3005] = -9'sd57;
	qsin_lut[3006] =  9'sd26;
	icos_lut[3006] = -9'sd64;
	qsin_lut[3007] =  9'sd13;
	icos_lut[3007] = -9'sd68;
	qsin_lut[3008] =  9'sd0;
	icos_lut[3008] = -9'sd67;
	qsin_lut[3009] = -9'sd13;
	icos_lut[3009] = -9'sd66;
	qsin_lut[3010] = -9'sd26;
	icos_lut[3010] = -9'sd62;
	qsin_lut[3011] = -9'sd37;
	icos_lut[3011] = -9'sd56;
	qsin_lut[3012] = -9'sd47;
	icos_lut[3012] = -9'sd47;
	qsin_lut[3013] = -9'sd56;
	icos_lut[3013] = -9'sd37;
	qsin_lut[3014] = -9'sd62;
	icos_lut[3014] = -9'sd26;
	qsin_lut[3015] = -9'sd66;
	icos_lut[3015] = -9'sd13;
	qsin_lut[3016] = -9'sd67;
	icos_lut[3016] = -9'sd0;
	qsin_lut[3017] = -9'sd66;
	icos_lut[3017] =  9'sd13;
	qsin_lut[3018] = -9'sd62;
	icos_lut[3018] =  9'sd26;
	qsin_lut[3019] = -9'sd56;
	icos_lut[3019] =  9'sd37;
	qsin_lut[3020] = -9'sd47;
	icos_lut[3020] =  9'sd47;
	qsin_lut[3021] = -9'sd37;
	icos_lut[3021] =  9'sd56;
	qsin_lut[3022] = -9'sd26;
	icos_lut[3022] =  9'sd62;
	qsin_lut[3023] = -9'sd13;
	icos_lut[3023] =  9'sd66;
	qsin_lut[3024] = -9'sd0;
	icos_lut[3024] =  9'sd67;
	qsin_lut[3025] =  9'sd13;
	icos_lut[3025] =  9'sd66;
	qsin_lut[3026] =  9'sd26;
	icos_lut[3026] =  9'sd62;
	qsin_lut[3027] =  9'sd37;
	icos_lut[3027] =  9'sd56;
	qsin_lut[3028] =  9'sd47;
	icos_lut[3028] =  9'sd47;
	qsin_lut[3029] =  9'sd56;
	icos_lut[3029] =  9'sd37;
	qsin_lut[3030] =  9'sd62;
	icos_lut[3030] =  9'sd26;
	qsin_lut[3031] =  9'sd66;
	icos_lut[3031] =  9'sd13;
	qsin_lut[3032] =  9'sd67;
	icos_lut[3032] =  9'sd0;
	qsin_lut[3033] =  9'sd66;
	icos_lut[3033] = -9'sd13;
	qsin_lut[3034] =  9'sd62;
	icos_lut[3034] = -9'sd26;
	qsin_lut[3035] =  9'sd56;
	icos_lut[3035] = -9'sd37;
	qsin_lut[3036] =  9'sd47;
	icos_lut[3036] = -9'sd47;
	qsin_lut[3037] =  9'sd37;
	icos_lut[3037] = -9'sd56;
	qsin_lut[3038] =  9'sd26;
	icos_lut[3038] = -9'sd62;
	qsin_lut[3039] =  9'sd13;
	icos_lut[3039] = -9'sd66;
	qsin_lut[3040] =  9'sd0;
	icos_lut[3040] = -9'sd65;
	qsin_lut[3041] = -9'sd13;
	icos_lut[3041] = -9'sd64;
	qsin_lut[3042] = -9'sd25;
	icos_lut[3042] = -9'sd60;
	qsin_lut[3043] = -9'sd36;
	icos_lut[3043] = -9'sd54;
	qsin_lut[3044] = -9'sd46;
	icos_lut[3044] = -9'sd46;
	qsin_lut[3045] = -9'sd54;
	icos_lut[3045] = -9'sd36;
	qsin_lut[3046] = -9'sd60;
	icos_lut[3046] = -9'sd25;
	qsin_lut[3047] = -9'sd64;
	icos_lut[3047] = -9'sd13;
	qsin_lut[3048] = -9'sd65;
	icos_lut[3048] = -9'sd0;
	qsin_lut[3049] = -9'sd64;
	icos_lut[3049] =  9'sd13;
	qsin_lut[3050] = -9'sd60;
	icos_lut[3050] =  9'sd25;
	qsin_lut[3051] = -9'sd54;
	icos_lut[3051] =  9'sd36;
	qsin_lut[3052] = -9'sd46;
	icos_lut[3052] =  9'sd46;
	qsin_lut[3053] = -9'sd36;
	icos_lut[3053] =  9'sd54;
	qsin_lut[3054] = -9'sd25;
	icos_lut[3054] =  9'sd60;
	qsin_lut[3055] = -9'sd13;
	icos_lut[3055] =  9'sd64;
	qsin_lut[3056] = -9'sd0;
	icos_lut[3056] =  9'sd65;
	qsin_lut[3057] =  9'sd13;
	icos_lut[3057] =  9'sd64;
	qsin_lut[3058] =  9'sd25;
	icos_lut[3058] =  9'sd60;
	qsin_lut[3059] =  9'sd36;
	icos_lut[3059] =  9'sd54;
	qsin_lut[3060] =  9'sd46;
	icos_lut[3060] =  9'sd46;
	qsin_lut[3061] =  9'sd54;
	icos_lut[3061] =  9'sd36;
	qsin_lut[3062] =  9'sd60;
	icos_lut[3062] =  9'sd25;
	qsin_lut[3063] =  9'sd64;
	icos_lut[3063] =  9'sd13;
	qsin_lut[3064] =  9'sd65;
	icos_lut[3064] =  9'sd0;
	qsin_lut[3065] =  9'sd64;
	icos_lut[3065] = -9'sd13;
	qsin_lut[3066] =  9'sd60;
	icos_lut[3066] = -9'sd25;
	qsin_lut[3067] =  9'sd54;
	icos_lut[3067] = -9'sd36;
	qsin_lut[3068] =  9'sd46;
	icos_lut[3068] = -9'sd46;
	qsin_lut[3069] =  9'sd36;
	icos_lut[3069] = -9'sd54;
	qsin_lut[3070] =  9'sd25;
	icos_lut[3070] = -9'sd60;
	qsin_lut[3071] =  9'sd13;
	icos_lut[3071] = -9'sd64;
	qsin_lut[3072] =  9'sd0;
	icos_lut[3072] = -9'sd63;
	qsin_lut[3073] = -9'sd12;
	icos_lut[3073] = -9'sd62;
	qsin_lut[3074] = -9'sd24;
	icos_lut[3074] = -9'sd58;
	qsin_lut[3075] = -9'sd35;
	icos_lut[3075] = -9'sd52;
	qsin_lut[3076] = -9'sd45;
	icos_lut[3076] = -9'sd45;
	qsin_lut[3077] = -9'sd52;
	icos_lut[3077] = -9'sd35;
	qsin_lut[3078] = -9'sd58;
	icos_lut[3078] = -9'sd24;
	qsin_lut[3079] = -9'sd62;
	icos_lut[3079] = -9'sd12;
	qsin_lut[3080] = -9'sd63;
	icos_lut[3080] = -9'sd0;
	qsin_lut[3081] = -9'sd62;
	icos_lut[3081] =  9'sd12;
	qsin_lut[3082] = -9'sd58;
	icos_lut[3082] =  9'sd24;
	qsin_lut[3083] = -9'sd52;
	icos_lut[3083] =  9'sd35;
	qsin_lut[3084] = -9'sd45;
	icos_lut[3084] =  9'sd45;
	qsin_lut[3085] = -9'sd35;
	icos_lut[3085] =  9'sd52;
	qsin_lut[3086] = -9'sd24;
	icos_lut[3086] =  9'sd58;
	qsin_lut[3087] = -9'sd12;
	icos_lut[3087] =  9'sd62;
	qsin_lut[3088] = -9'sd0;
	icos_lut[3088] =  9'sd63;
	qsin_lut[3089] =  9'sd12;
	icos_lut[3089] =  9'sd62;
	qsin_lut[3090] =  9'sd24;
	icos_lut[3090] =  9'sd58;
	qsin_lut[3091] =  9'sd35;
	icos_lut[3091] =  9'sd52;
	qsin_lut[3092] =  9'sd45;
	icos_lut[3092] =  9'sd45;
	qsin_lut[3093] =  9'sd52;
	icos_lut[3093] =  9'sd35;
	qsin_lut[3094] =  9'sd58;
	icos_lut[3094] =  9'sd24;
	qsin_lut[3095] =  9'sd62;
	icos_lut[3095] =  9'sd12;
	qsin_lut[3096] =  9'sd63;
	icos_lut[3096] =  9'sd0;
	qsin_lut[3097] =  9'sd62;
	icos_lut[3097] = -9'sd12;
	qsin_lut[3098] =  9'sd58;
	icos_lut[3098] = -9'sd24;
	qsin_lut[3099] =  9'sd52;
	icos_lut[3099] = -9'sd35;
	qsin_lut[3100] =  9'sd45;
	icos_lut[3100] = -9'sd45;
	qsin_lut[3101] =  9'sd35;
	icos_lut[3101] = -9'sd52;
	qsin_lut[3102] =  9'sd24;
	icos_lut[3102] = -9'sd58;
	qsin_lut[3103] =  9'sd12;
	icos_lut[3103] = -9'sd62;
	qsin_lut[3104] =  9'sd0;
	icos_lut[3104] = -9'sd61;
	qsin_lut[3105] = -9'sd12;
	icos_lut[3105] = -9'sd60;
	qsin_lut[3106] = -9'sd23;
	icos_lut[3106] = -9'sd56;
	qsin_lut[3107] = -9'sd34;
	icos_lut[3107] = -9'sd51;
	qsin_lut[3108] = -9'sd43;
	icos_lut[3108] = -9'sd43;
	qsin_lut[3109] = -9'sd51;
	icos_lut[3109] = -9'sd34;
	qsin_lut[3110] = -9'sd56;
	icos_lut[3110] = -9'sd23;
	qsin_lut[3111] = -9'sd60;
	icos_lut[3111] = -9'sd12;
	qsin_lut[3112] = -9'sd61;
	icos_lut[3112] = -9'sd0;
	qsin_lut[3113] = -9'sd60;
	icos_lut[3113] =  9'sd12;
	qsin_lut[3114] = -9'sd56;
	icos_lut[3114] =  9'sd23;
	qsin_lut[3115] = -9'sd51;
	icos_lut[3115] =  9'sd34;
	qsin_lut[3116] = -9'sd43;
	icos_lut[3116] =  9'sd43;
	qsin_lut[3117] = -9'sd34;
	icos_lut[3117] =  9'sd51;
	qsin_lut[3118] = -9'sd23;
	icos_lut[3118] =  9'sd56;
	qsin_lut[3119] = -9'sd12;
	icos_lut[3119] =  9'sd60;
	qsin_lut[3120] = -9'sd0;
	icos_lut[3120] =  9'sd61;
	qsin_lut[3121] =  9'sd12;
	icos_lut[3121] =  9'sd60;
	qsin_lut[3122] =  9'sd23;
	icos_lut[3122] =  9'sd56;
	qsin_lut[3123] =  9'sd34;
	icos_lut[3123] =  9'sd51;
	qsin_lut[3124] =  9'sd43;
	icos_lut[3124] =  9'sd43;
	qsin_lut[3125] =  9'sd51;
	icos_lut[3125] =  9'sd34;
	qsin_lut[3126] =  9'sd56;
	icos_lut[3126] =  9'sd23;
	qsin_lut[3127] =  9'sd60;
	icos_lut[3127] =  9'sd12;
	qsin_lut[3128] =  9'sd61;
	icos_lut[3128] =  9'sd0;
	qsin_lut[3129] =  9'sd60;
	icos_lut[3129] = -9'sd12;
	qsin_lut[3130] =  9'sd56;
	icos_lut[3130] = -9'sd23;
	qsin_lut[3131] =  9'sd51;
	icos_lut[3131] = -9'sd34;
	qsin_lut[3132] =  9'sd43;
	icos_lut[3132] = -9'sd43;
	qsin_lut[3133] =  9'sd34;
	icos_lut[3133] = -9'sd51;
	qsin_lut[3134] =  9'sd23;
	icos_lut[3134] = -9'sd56;
	qsin_lut[3135] =  9'sd12;
	icos_lut[3135] = -9'sd60;
	qsin_lut[3136] =  9'sd0;
	icos_lut[3136] = -9'sd59;
	qsin_lut[3137] = -9'sd12;
	icos_lut[3137] = -9'sd58;
	qsin_lut[3138] = -9'sd23;
	icos_lut[3138] = -9'sd55;
	qsin_lut[3139] = -9'sd33;
	icos_lut[3139] = -9'sd49;
	qsin_lut[3140] = -9'sd42;
	icos_lut[3140] = -9'sd42;
	qsin_lut[3141] = -9'sd49;
	icos_lut[3141] = -9'sd33;
	qsin_lut[3142] = -9'sd55;
	icos_lut[3142] = -9'sd23;
	qsin_lut[3143] = -9'sd58;
	icos_lut[3143] = -9'sd12;
	qsin_lut[3144] = -9'sd59;
	icos_lut[3144] = -9'sd0;
	qsin_lut[3145] = -9'sd58;
	icos_lut[3145] =  9'sd12;
	qsin_lut[3146] = -9'sd55;
	icos_lut[3146] =  9'sd23;
	qsin_lut[3147] = -9'sd49;
	icos_lut[3147] =  9'sd33;
	qsin_lut[3148] = -9'sd42;
	icos_lut[3148] =  9'sd42;
	qsin_lut[3149] = -9'sd33;
	icos_lut[3149] =  9'sd49;
	qsin_lut[3150] = -9'sd23;
	icos_lut[3150] =  9'sd55;
	qsin_lut[3151] = -9'sd12;
	icos_lut[3151] =  9'sd58;
	qsin_lut[3152] = -9'sd0;
	icos_lut[3152] =  9'sd59;
	qsin_lut[3153] =  9'sd12;
	icos_lut[3153] =  9'sd58;
	qsin_lut[3154] =  9'sd23;
	icos_lut[3154] =  9'sd55;
	qsin_lut[3155] =  9'sd33;
	icos_lut[3155] =  9'sd49;
	qsin_lut[3156] =  9'sd42;
	icos_lut[3156] =  9'sd42;
	qsin_lut[3157] =  9'sd49;
	icos_lut[3157] =  9'sd33;
	qsin_lut[3158] =  9'sd55;
	icos_lut[3158] =  9'sd23;
	qsin_lut[3159] =  9'sd58;
	icos_lut[3159] =  9'sd12;
	qsin_lut[3160] =  9'sd59;
	icos_lut[3160] =  9'sd0;
	qsin_lut[3161] =  9'sd58;
	icos_lut[3161] = -9'sd12;
	qsin_lut[3162] =  9'sd55;
	icos_lut[3162] = -9'sd23;
	qsin_lut[3163] =  9'sd49;
	icos_lut[3163] = -9'sd33;
	qsin_lut[3164] =  9'sd42;
	icos_lut[3164] = -9'sd42;
	qsin_lut[3165] =  9'sd33;
	icos_lut[3165] = -9'sd49;
	qsin_lut[3166] =  9'sd23;
	icos_lut[3166] = -9'sd55;
	qsin_lut[3167] =  9'sd12;
	icos_lut[3167] = -9'sd58;
	qsin_lut[3168] =  9'sd0;
	icos_lut[3168] = -9'sd57;
	qsin_lut[3169] = -9'sd11;
	icos_lut[3169] = -9'sd56;
	qsin_lut[3170] = -9'sd22;
	icos_lut[3170] = -9'sd53;
	qsin_lut[3171] = -9'sd32;
	icos_lut[3171] = -9'sd47;
	qsin_lut[3172] = -9'sd40;
	icos_lut[3172] = -9'sd40;
	qsin_lut[3173] = -9'sd47;
	icos_lut[3173] = -9'sd32;
	qsin_lut[3174] = -9'sd53;
	icos_lut[3174] = -9'sd22;
	qsin_lut[3175] = -9'sd56;
	icos_lut[3175] = -9'sd11;
	qsin_lut[3176] = -9'sd57;
	icos_lut[3176] = -9'sd0;
	qsin_lut[3177] = -9'sd56;
	icos_lut[3177] =  9'sd11;
	qsin_lut[3178] = -9'sd53;
	icos_lut[3178] =  9'sd22;
	qsin_lut[3179] = -9'sd47;
	icos_lut[3179] =  9'sd32;
	qsin_lut[3180] = -9'sd40;
	icos_lut[3180] =  9'sd40;
	qsin_lut[3181] = -9'sd32;
	icos_lut[3181] =  9'sd47;
	qsin_lut[3182] = -9'sd22;
	icos_lut[3182] =  9'sd53;
	qsin_lut[3183] = -9'sd11;
	icos_lut[3183] =  9'sd56;
	qsin_lut[3184] = -9'sd0;
	icos_lut[3184] =  9'sd57;
	qsin_lut[3185] =  9'sd11;
	icos_lut[3185] =  9'sd56;
	qsin_lut[3186] =  9'sd22;
	icos_lut[3186] =  9'sd53;
	qsin_lut[3187] =  9'sd32;
	icos_lut[3187] =  9'sd47;
	qsin_lut[3188] =  9'sd40;
	icos_lut[3188] =  9'sd40;
	qsin_lut[3189] =  9'sd47;
	icos_lut[3189] =  9'sd32;
	qsin_lut[3190] =  9'sd53;
	icos_lut[3190] =  9'sd22;
	qsin_lut[3191] =  9'sd56;
	icos_lut[3191] =  9'sd11;
	qsin_lut[3192] =  9'sd57;
	icos_lut[3192] =  9'sd0;
	qsin_lut[3193] =  9'sd56;
	icos_lut[3193] = -9'sd11;
	qsin_lut[3194] =  9'sd53;
	icos_lut[3194] = -9'sd22;
	qsin_lut[3195] =  9'sd47;
	icos_lut[3195] = -9'sd32;
	qsin_lut[3196] =  9'sd40;
	icos_lut[3196] = -9'sd40;
	qsin_lut[3197] =  9'sd32;
	icos_lut[3197] = -9'sd47;
	qsin_lut[3198] =  9'sd22;
	icos_lut[3198] = -9'sd53;
	qsin_lut[3199] =  9'sd11;
	icos_lut[3199] = -9'sd56;
	qsin_lut[3200] =  9'sd0;
	icos_lut[3200] = -9'sd55;
	qsin_lut[3201] = -9'sd11;
	icos_lut[3201] = -9'sd54;
	qsin_lut[3202] = -9'sd21;
	icos_lut[3202] = -9'sd51;
	qsin_lut[3203] = -9'sd31;
	icos_lut[3203] = -9'sd46;
	qsin_lut[3204] = -9'sd39;
	icos_lut[3204] = -9'sd39;
	qsin_lut[3205] = -9'sd46;
	icos_lut[3205] = -9'sd31;
	qsin_lut[3206] = -9'sd51;
	icos_lut[3206] = -9'sd21;
	qsin_lut[3207] = -9'sd54;
	icos_lut[3207] = -9'sd11;
	qsin_lut[3208] = -9'sd55;
	icos_lut[3208] = -9'sd0;
	qsin_lut[3209] = -9'sd54;
	icos_lut[3209] =  9'sd11;
	qsin_lut[3210] = -9'sd51;
	icos_lut[3210] =  9'sd21;
	qsin_lut[3211] = -9'sd46;
	icos_lut[3211] =  9'sd31;
	qsin_lut[3212] = -9'sd39;
	icos_lut[3212] =  9'sd39;
	qsin_lut[3213] = -9'sd31;
	icos_lut[3213] =  9'sd46;
	qsin_lut[3214] = -9'sd21;
	icos_lut[3214] =  9'sd51;
	qsin_lut[3215] = -9'sd11;
	icos_lut[3215] =  9'sd54;
	qsin_lut[3216] = -9'sd0;
	icos_lut[3216] =  9'sd55;
	qsin_lut[3217] =  9'sd11;
	icos_lut[3217] =  9'sd54;
	qsin_lut[3218] =  9'sd21;
	icos_lut[3218] =  9'sd51;
	qsin_lut[3219] =  9'sd31;
	icos_lut[3219] =  9'sd46;
	qsin_lut[3220] =  9'sd39;
	icos_lut[3220] =  9'sd39;
	qsin_lut[3221] =  9'sd46;
	icos_lut[3221] =  9'sd31;
	qsin_lut[3222] =  9'sd51;
	icos_lut[3222] =  9'sd21;
	qsin_lut[3223] =  9'sd54;
	icos_lut[3223] =  9'sd11;
	qsin_lut[3224] =  9'sd55;
	icos_lut[3224] =  9'sd0;
	qsin_lut[3225] =  9'sd54;
	icos_lut[3225] = -9'sd11;
	qsin_lut[3226] =  9'sd51;
	icos_lut[3226] = -9'sd21;
	qsin_lut[3227] =  9'sd46;
	icos_lut[3227] = -9'sd31;
	qsin_lut[3228] =  9'sd39;
	icos_lut[3228] = -9'sd39;
	qsin_lut[3229] =  9'sd31;
	icos_lut[3229] = -9'sd46;
	qsin_lut[3230] =  9'sd21;
	icos_lut[3230] = -9'sd51;
	qsin_lut[3231] =  9'sd11;
	icos_lut[3231] = -9'sd54;
	qsin_lut[3232] =  9'sd0;
	icos_lut[3232] = -9'sd53;
	qsin_lut[3233] = -9'sd10;
	icos_lut[3233] = -9'sd52;
	qsin_lut[3234] = -9'sd20;
	icos_lut[3234] = -9'sd49;
	qsin_lut[3235] = -9'sd29;
	icos_lut[3235] = -9'sd44;
	qsin_lut[3236] = -9'sd37;
	icos_lut[3236] = -9'sd37;
	qsin_lut[3237] = -9'sd44;
	icos_lut[3237] = -9'sd29;
	qsin_lut[3238] = -9'sd49;
	icos_lut[3238] = -9'sd20;
	qsin_lut[3239] = -9'sd52;
	icos_lut[3239] = -9'sd10;
	qsin_lut[3240] = -9'sd53;
	icos_lut[3240] = -9'sd0;
	qsin_lut[3241] = -9'sd52;
	icos_lut[3241] =  9'sd10;
	qsin_lut[3242] = -9'sd49;
	icos_lut[3242] =  9'sd20;
	qsin_lut[3243] = -9'sd44;
	icos_lut[3243] =  9'sd29;
	qsin_lut[3244] = -9'sd37;
	icos_lut[3244] =  9'sd37;
	qsin_lut[3245] = -9'sd29;
	icos_lut[3245] =  9'sd44;
	qsin_lut[3246] = -9'sd20;
	icos_lut[3246] =  9'sd49;
	qsin_lut[3247] = -9'sd10;
	icos_lut[3247] =  9'sd52;
	qsin_lut[3248] = -9'sd0;
	icos_lut[3248] =  9'sd53;
	qsin_lut[3249] =  9'sd10;
	icos_lut[3249] =  9'sd52;
	qsin_lut[3250] =  9'sd20;
	icos_lut[3250] =  9'sd49;
	qsin_lut[3251] =  9'sd29;
	icos_lut[3251] =  9'sd44;
	qsin_lut[3252] =  9'sd37;
	icos_lut[3252] =  9'sd37;
	qsin_lut[3253] =  9'sd44;
	icos_lut[3253] =  9'sd29;
	qsin_lut[3254] =  9'sd49;
	icos_lut[3254] =  9'sd20;
	qsin_lut[3255] =  9'sd52;
	icos_lut[3255] =  9'sd10;
	qsin_lut[3256] =  9'sd53;
	icos_lut[3256] =  9'sd0;
	qsin_lut[3257] =  9'sd52;
	icos_lut[3257] = -9'sd10;
	qsin_lut[3258] =  9'sd49;
	icos_lut[3258] = -9'sd20;
	qsin_lut[3259] =  9'sd44;
	icos_lut[3259] = -9'sd29;
	qsin_lut[3260] =  9'sd37;
	icos_lut[3260] = -9'sd37;
	qsin_lut[3261] =  9'sd29;
	icos_lut[3261] = -9'sd44;
	qsin_lut[3262] =  9'sd20;
	icos_lut[3262] = -9'sd49;
	qsin_lut[3263] =  9'sd10;
	icos_lut[3263] = -9'sd52;
	qsin_lut[3264] =  9'sd0;
	icos_lut[3264] = -9'sd51;
	qsin_lut[3265] = -9'sd10;
	icos_lut[3265] = -9'sd50;
	qsin_lut[3266] = -9'sd20;
	icos_lut[3266] = -9'sd47;
	qsin_lut[3267] = -9'sd28;
	icos_lut[3267] = -9'sd42;
	qsin_lut[3268] = -9'sd36;
	icos_lut[3268] = -9'sd36;
	qsin_lut[3269] = -9'sd42;
	icos_lut[3269] = -9'sd28;
	qsin_lut[3270] = -9'sd47;
	icos_lut[3270] = -9'sd20;
	qsin_lut[3271] = -9'sd50;
	icos_lut[3271] = -9'sd10;
	qsin_lut[3272] = -9'sd51;
	icos_lut[3272] = -9'sd0;
	qsin_lut[3273] = -9'sd50;
	icos_lut[3273] =  9'sd10;
	qsin_lut[3274] = -9'sd47;
	icos_lut[3274] =  9'sd20;
	qsin_lut[3275] = -9'sd42;
	icos_lut[3275] =  9'sd28;
	qsin_lut[3276] = -9'sd36;
	icos_lut[3276] =  9'sd36;
	qsin_lut[3277] = -9'sd28;
	icos_lut[3277] =  9'sd42;
	qsin_lut[3278] = -9'sd20;
	icos_lut[3278] =  9'sd47;
	qsin_lut[3279] = -9'sd10;
	icos_lut[3279] =  9'sd50;
	qsin_lut[3280] = -9'sd0;
	icos_lut[3280] =  9'sd51;
	qsin_lut[3281] =  9'sd10;
	icos_lut[3281] =  9'sd50;
	qsin_lut[3282] =  9'sd20;
	icos_lut[3282] =  9'sd47;
	qsin_lut[3283] =  9'sd28;
	icos_lut[3283] =  9'sd42;
	qsin_lut[3284] =  9'sd36;
	icos_lut[3284] =  9'sd36;
	qsin_lut[3285] =  9'sd42;
	icos_lut[3285] =  9'sd28;
	qsin_lut[3286] =  9'sd47;
	icos_lut[3286] =  9'sd20;
	qsin_lut[3287] =  9'sd50;
	icos_lut[3287] =  9'sd10;
	qsin_lut[3288] =  9'sd51;
	icos_lut[3288] =  9'sd0;
	qsin_lut[3289] =  9'sd50;
	icos_lut[3289] = -9'sd10;
	qsin_lut[3290] =  9'sd47;
	icos_lut[3290] = -9'sd20;
	qsin_lut[3291] =  9'sd42;
	icos_lut[3291] = -9'sd28;
	qsin_lut[3292] =  9'sd36;
	icos_lut[3292] = -9'sd36;
	qsin_lut[3293] =  9'sd28;
	icos_lut[3293] = -9'sd42;
	qsin_lut[3294] =  9'sd20;
	icos_lut[3294] = -9'sd47;
	qsin_lut[3295] =  9'sd10;
	icos_lut[3295] = -9'sd50;
	qsin_lut[3296] =  9'sd0;
	icos_lut[3296] = -9'sd49;
	qsin_lut[3297] = -9'sd10;
	icos_lut[3297] = -9'sd48;
	qsin_lut[3298] = -9'sd19;
	icos_lut[3298] = -9'sd45;
	qsin_lut[3299] = -9'sd27;
	icos_lut[3299] = -9'sd41;
	qsin_lut[3300] = -9'sd35;
	icos_lut[3300] = -9'sd35;
	qsin_lut[3301] = -9'sd41;
	icos_lut[3301] = -9'sd27;
	qsin_lut[3302] = -9'sd45;
	icos_lut[3302] = -9'sd19;
	qsin_lut[3303] = -9'sd48;
	icos_lut[3303] = -9'sd10;
	qsin_lut[3304] = -9'sd49;
	icos_lut[3304] = -9'sd0;
	qsin_lut[3305] = -9'sd48;
	icos_lut[3305] =  9'sd10;
	qsin_lut[3306] = -9'sd45;
	icos_lut[3306] =  9'sd19;
	qsin_lut[3307] = -9'sd41;
	icos_lut[3307] =  9'sd27;
	qsin_lut[3308] = -9'sd35;
	icos_lut[3308] =  9'sd35;
	qsin_lut[3309] = -9'sd27;
	icos_lut[3309] =  9'sd41;
	qsin_lut[3310] = -9'sd19;
	icos_lut[3310] =  9'sd45;
	qsin_lut[3311] = -9'sd10;
	icos_lut[3311] =  9'sd48;
	qsin_lut[3312] = -9'sd0;
	icos_lut[3312] =  9'sd49;
	qsin_lut[3313] =  9'sd10;
	icos_lut[3313] =  9'sd48;
	qsin_lut[3314] =  9'sd19;
	icos_lut[3314] =  9'sd45;
	qsin_lut[3315] =  9'sd27;
	icos_lut[3315] =  9'sd41;
	qsin_lut[3316] =  9'sd35;
	icos_lut[3316] =  9'sd35;
	qsin_lut[3317] =  9'sd41;
	icos_lut[3317] =  9'sd27;
	qsin_lut[3318] =  9'sd45;
	icos_lut[3318] =  9'sd19;
	qsin_lut[3319] =  9'sd48;
	icos_lut[3319] =  9'sd10;
	qsin_lut[3320] =  9'sd49;
	icos_lut[3320] =  9'sd0;
	qsin_lut[3321] =  9'sd48;
	icos_lut[3321] = -9'sd10;
	qsin_lut[3322] =  9'sd45;
	icos_lut[3322] = -9'sd19;
	qsin_lut[3323] =  9'sd41;
	icos_lut[3323] = -9'sd27;
	qsin_lut[3324] =  9'sd35;
	icos_lut[3324] = -9'sd35;
	qsin_lut[3325] =  9'sd27;
	icos_lut[3325] = -9'sd41;
	qsin_lut[3326] =  9'sd19;
	icos_lut[3326] = -9'sd45;
	qsin_lut[3327] =  9'sd10;
	icos_lut[3327] = -9'sd48;
	qsin_lut[3328] =  9'sd0;
	icos_lut[3328] = -9'sd47;
	qsin_lut[3329] = -9'sd9;
	icos_lut[3329] = -9'sd46;
	qsin_lut[3330] = -9'sd18;
	icos_lut[3330] = -9'sd43;
	qsin_lut[3331] = -9'sd26;
	icos_lut[3331] = -9'sd39;
	qsin_lut[3332] = -9'sd33;
	icos_lut[3332] = -9'sd33;
	qsin_lut[3333] = -9'sd39;
	icos_lut[3333] = -9'sd26;
	qsin_lut[3334] = -9'sd43;
	icos_lut[3334] = -9'sd18;
	qsin_lut[3335] = -9'sd46;
	icos_lut[3335] = -9'sd9;
	qsin_lut[3336] = -9'sd47;
	icos_lut[3336] = -9'sd0;
	qsin_lut[3337] = -9'sd46;
	icos_lut[3337] =  9'sd9;
	qsin_lut[3338] = -9'sd43;
	icos_lut[3338] =  9'sd18;
	qsin_lut[3339] = -9'sd39;
	icos_lut[3339] =  9'sd26;
	qsin_lut[3340] = -9'sd33;
	icos_lut[3340] =  9'sd33;
	qsin_lut[3341] = -9'sd26;
	icos_lut[3341] =  9'sd39;
	qsin_lut[3342] = -9'sd18;
	icos_lut[3342] =  9'sd43;
	qsin_lut[3343] = -9'sd9;
	icos_lut[3343] =  9'sd46;
	qsin_lut[3344] = -9'sd0;
	icos_lut[3344] =  9'sd47;
	qsin_lut[3345] =  9'sd9;
	icos_lut[3345] =  9'sd46;
	qsin_lut[3346] =  9'sd18;
	icos_lut[3346] =  9'sd43;
	qsin_lut[3347] =  9'sd26;
	icos_lut[3347] =  9'sd39;
	qsin_lut[3348] =  9'sd33;
	icos_lut[3348] =  9'sd33;
	qsin_lut[3349] =  9'sd39;
	icos_lut[3349] =  9'sd26;
	qsin_lut[3350] =  9'sd43;
	icos_lut[3350] =  9'sd18;
	qsin_lut[3351] =  9'sd46;
	icos_lut[3351] =  9'sd9;
	qsin_lut[3352] =  9'sd47;
	icos_lut[3352] =  9'sd0;
	qsin_lut[3353] =  9'sd46;
	icos_lut[3353] = -9'sd9;
	qsin_lut[3354] =  9'sd43;
	icos_lut[3354] = -9'sd18;
	qsin_lut[3355] =  9'sd39;
	icos_lut[3355] = -9'sd26;
	qsin_lut[3356] =  9'sd33;
	icos_lut[3356] = -9'sd33;
	qsin_lut[3357] =  9'sd26;
	icos_lut[3357] = -9'sd39;
	qsin_lut[3358] =  9'sd18;
	icos_lut[3358] = -9'sd43;
	qsin_lut[3359] =  9'sd9;
	icos_lut[3359] = -9'sd46;
	qsin_lut[3360] =  9'sd0;
	icos_lut[3360] = -9'sd45;
	qsin_lut[3361] = -9'sd9;
	icos_lut[3361] = -9'sd44;
	qsin_lut[3362] = -9'sd17;
	icos_lut[3362] = -9'sd42;
	qsin_lut[3363] = -9'sd25;
	icos_lut[3363] = -9'sd37;
	qsin_lut[3364] = -9'sd32;
	icos_lut[3364] = -9'sd32;
	qsin_lut[3365] = -9'sd37;
	icos_lut[3365] = -9'sd25;
	qsin_lut[3366] = -9'sd42;
	icos_lut[3366] = -9'sd17;
	qsin_lut[3367] = -9'sd44;
	icos_lut[3367] = -9'sd9;
	qsin_lut[3368] = -9'sd45;
	icos_lut[3368] = -9'sd0;
	qsin_lut[3369] = -9'sd44;
	icos_lut[3369] =  9'sd9;
	qsin_lut[3370] = -9'sd42;
	icos_lut[3370] =  9'sd17;
	qsin_lut[3371] = -9'sd37;
	icos_lut[3371] =  9'sd25;
	qsin_lut[3372] = -9'sd32;
	icos_lut[3372] =  9'sd32;
	qsin_lut[3373] = -9'sd25;
	icos_lut[3373] =  9'sd37;
	qsin_lut[3374] = -9'sd17;
	icos_lut[3374] =  9'sd42;
	qsin_lut[3375] = -9'sd9;
	icos_lut[3375] =  9'sd44;
	qsin_lut[3376] = -9'sd0;
	icos_lut[3376] =  9'sd45;
	qsin_lut[3377] =  9'sd9;
	icos_lut[3377] =  9'sd44;
	qsin_lut[3378] =  9'sd17;
	icos_lut[3378] =  9'sd42;
	qsin_lut[3379] =  9'sd25;
	icos_lut[3379] =  9'sd37;
	qsin_lut[3380] =  9'sd32;
	icos_lut[3380] =  9'sd32;
	qsin_lut[3381] =  9'sd37;
	icos_lut[3381] =  9'sd25;
	qsin_lut[3382] =  9'sd42;
	icos_lut[3382] =  9'sd17;
	qsin_lut[3383] =  9'sd44;
	icos_lut[3383] =  9'sd9;
	qsin_lut[3384] =  9'sd45;
	icos_lut[3384] =  9'sd0;
	qsin_lut[3385] =  9'sd44;
	icos_lut[3385] = -9'sd9;
	qsin_lut[3386] =  9'sd42;
	icos_lut[3386] = -9'sd17;
	qsin_lut[3387] =  9'sd37;
	icos_lut[3387] = -9'sd25;
	qsin_lut[3388] =  9'sd32;
	icos_lut[3388] = -9'sd32;
	qsin_lut[3389] =  9'sd25;
	icos_lut[3389] = -9'sd37;
	qsin_lut[3390] =  9'sd17;
	icos_lut[3390] = -9'sd42;
	qsin_lut[3391] =  9'sd9;
	icos_lut[3391] = -9'sd44;
	qsin_lut[3392] =  9'sd0;
	icos_lut[3392] = -9'sd43;
	qsin_lut[3393] = -9'sd8;
	icos_lut[3393] = -9'sd42;
	qsin_lut[3394] = -9'sd16;
	icos_lut[3394] = -9'sd40;
	qsin_lut[3395] = -9'sd24;
	icos_lut[3395] = -9'sd36;
	qsin_lut[3396] = -9'sd30;
	icos_lut[3396] = -9'sd30;
	qsin_lut[3397] = -9'sd36;
	icos_lut[3397] = -9'sd24;
	qsin_lut[3398] = -9'sd40;
	icos_lut[3398] = -9'sd16;
	qsin_lut[3399] = -9'sd42;
	icos_lut[3399] = -9'sd8;
	qsin_lut[3400] = -9'sd43;
	icos_lut[3400] = -9'sd0;
	qsin_lut[3401] = -9'sd42;
	icos_lut[3401] =  9'sd8;
	qsin_lut[3402] = -9'sd40;
	icos_lut[3402] =  9'sd16;
	qsin_lut[3403] = -9'sd36;
	icos_lut[3403] =  9'sd24;
	qsin_lut[3404] = -9'sd30;
	icos_lut[3404] =  9'sd30;
	qsin_lut[3405] = -9'sd24;
	icos_lut[3405] =  9'sd36;
	qsin_lut[3406] = -9'sd16;
	icos_lut[3406] =  9'sd40;
	qsin_lut[3407] = -9'sd8;
	icos_lut[3407] =  9'sd42;
	qsin_lut[3408] = -9'sd0;
	icos_lut[3408] =  9'sd43;
	qsin_lut[3409] =  9'sd8;
	icos_lut[3409] =  9'sd42;
	qsin_lut[3410] =  9'sd16;
	icos_lut[3410] =  9'sd40;
	qsin_lut[3411] =  9'sd24;
	icos_lut[3411] =  9'sd36;
	qsin_lut[3412] =  9'sd30;
	icos_lut[3412] =  9'sd30;
	qsin_lut[3413] =  9'sd36;
	icos_lut[3413] =  9'sd24;
	qsin_lut[3414] =  9'sd40;
	icos_lut[3414] =  9'sd16;
	qsin_lut[3415] =  9'sd42;
	icos_lut[3415] =  9'sd8;
	qsin_lut[3416] =  9'sd43;
	icos_lut[3416] =  9'sd0;
	qsin_lut[3417] =  9'sd42;
	icos_lut[3417] = -9'sd8;
	qsin_lut[3418] =  9'sd40;
	icos_lut[3418] = -9'sd16;
	qsin_lut[3419] =  9'sd36;
	icos_lut[3419] = -9'sd24;
	qsin_lut[3420] =  9'sd30;
	icos_lut[3420] = -9'sd30;
	qsin_lut[3421] =  9'sd24;
	icos_lut[3421] = -9'sd36;
	qsin_lut[3422] =  9'sd16;
	icos_lut[3422] = -9'sd40;
	qsin_lut[3423] =  9'sd8;
	icos_lut[3423] = -9'sd42;
	qsin_lut[3424] =  9'sd0;
	icos_lut[3424] = -9'sd41;
	qsin_lut[3425] = -9'sd8;
	icos_lut[3425] = -9'sd40;
	qsin_lut[3426] = -9'sd16;
	icos_lut[3426] = -9'sd38;
	qsin_lut[3427] = -9'sd23;
	icos_lut[3427] = -9'sd34;
	qsin_lut[3428] = -9'sd29;
	icos_lut[3428] = -9'sd29;
	qsin_lut[3429] = -9'sd34;
	icos_lut[3429] = -9'sd23;
	qsin_lut[3430] = -9'sd38;
	icos_lut[3430] = -9'sd16;
	qsin_lut[3431] = -9'sd40;
	icos_lut[3431] = -9'sd8;
	qsin_lut[3432] = -9'sd41;
	icos_lut[3432] = -9'sd0;
	qsin_lut[3433] = -9'sd40;
	icos_lut[3433] =  9'sd8;
	qsin_lut[3434] = -9'sd38;
	icos_lut[3434] =  9'sd16;
	qsin_lut[3435] = -9'sd34;
	icos_lut[3435] =  9'sd23;
	qsin_lut[3436] = -9'sd29;
	icos_lut[3436] =  9'sd29;
	qsin_lut[3437] = -9'sd23;
	icos_lut[3437] =  9'sd34;
	qsin_lut[3438] = -9'sd16;
	icos_lut[3438] =  9'sd38;
	qsin_lut[3439] = -9'sd8;
	icos_lut[3439] =  9'sd40;
	qsin_lut[3440] = -9'sd0;
	icos_lut[3440] =  9'sd41;
	qsin_lut[3441] =  9'sd8;
	icos_lut[3441] =  9'sd40;
	qsin_lut[3442] =  9'sd16;
	icos_lut[3442] =  9'sd38;
	qsin_lut[3443] =  9'sd23;
	icos_lut[3443] =  9'sd34;
	qsin_lut[3444] =  9'sd29;
	icos_lut[3444] =  9'sd29;
	qsin_lut[3445] =  9'sd34;
	icos_lut[3445] =  9'sd23;
	qsin_lut[3446] =  9'sd38;
	icos_lut[3446] =  9'sd16;
	qsin_lut[3447] =  9'sd40;
	icos_lut[3447] =  9'sd8;
	qsin_lut[3448] =  9'sd41;
	icos_lut[3448] =  9'sd0;
	qsin_lut[3449] =  9'sd40;
	icos_lut[3449] = -9'sd8;
	qsin_lut[3450] =  9'sd38;
	icos_lut[3450] = -9'sd16;
	qsin_lut[3451] =  9'sd34;
	icos_lut[3451] = -9'sd23;
	qsin_lut[3452] =  9'sd29;
	icos_lut[3452] = -9'sd29;
	qsin_lut[3453] =  9'sd23;
	icos_lut[3453] = -9'sd34;
	qsin_lut[3454] =  9'sd16;
	icos_lut[3454] = -9'sd38;
	qsin_lut[3455] =  9'sd8;
	icos_lut[3455] = -9'sd40;
	qsin_lut[3456] =  9'sd0;
	icos_lut[3456] = -9'sd39;
	qsin_lut[3457] = -9'sd8;
	icos_lut[3457] = -9'sd38;
	qsin_lut[3458] = -9'sd15;
	icos_lut[3458] = -9'sd36;
	qsin_lut[3459] = -9'sd22;
	icos_lut[3459] = -9'sd32;
	qsin_lut[3460] = -9'sd28;
	icos_lut[3460] = -9'sd28;
	qsin_lut[3461] = -9'sd32;
	icos_lut[3461] = -9'sd22;
	qsin_lut[3462] = -9'sd36;
	icos_lut[3462] = -9'sd15;
	qsin_lut[3463] = -9'sd38;
	icos_lut[3463] = -9'sd8;
	qsin_lut[3464] = -9'sd39;
	icos_lut[3464] = -9'sd0;
	qsin_lut[3465] = -9'sd38;
	icos_lut[3465] =  9'sd8;
	qsin_lut[3466] = -9'sd36;
	icos_lut[3466] =  9'sd15;
	qsin_lut[3467] = -9'sd32;
	icos_lut[3467] =  9'sd22;
	qsin_lut[3468] = -9'sd28;
	icos_lut[3468] =  9'sd28;
	qsin_lut[3469] = -9'sd22;
	icos_lut[3469] =  9'sd32;
	qsin_lut[3470] = -9'sd15;
	icos_lut[3470] =  9'sd36;
	qsin_lut[3471] = -9'sd8;
	icos_lut[3471] =  9'sd38;
	qsin_lut[3472] = -9'sd0;
	icos_lut[3472] =  9'sd39;
	qsin_lut[3473] =  9'sd8;
	icos_lut[3473] =  9'sd38;
	qsin_lut[3474] =  9'sd15;
	icos_lut[3474] =  9'sd36;
	qsin_lut[3475] =  9'sd22;
	icos_lut[3475] =  9'sd32;
	qsin_lut[3476] =  9'sd28;
	icos_lut[3476] =  9'sd28;
	qsin_lut[3477] =  9'sd32;
	icos_lut[3477] =  9'sd22;
	qsin_lut[3478] =  9'sd36;
	icos_lut[3478] =  9'sd15;
	qsin_lut[3479] =  9'sd38;
	icos_lut[3479] =  9'sd8;
	qsin_lut[3480] =  9'sd39;
	icos_lut[3480] =  9'sd0;
	qsin_lut[3481] =  9'sd38;
	icos_lut[3481] = -9'sd8;
	qsin_lut[3482] =  9'sd36;
	icos_lut[3482] = -9'sd15;
	qsin_lut[3483] =  9'sd32;
	icos_lut[3483] = -9'sd22;
	qsin_lut[3484] =  9'sd28;
	icos_lut[3484] = -9'sd28;
	qsin_lut[3485] =  9'sd22;
	icos_lut[3485] = -9'sd32;
	qsin_lut[3486] =  9'sd15;
	icos_lut[3486] = -9'sd36;
	qsin_lut[3487] =  9'sd8;
	icos_lut[3487] = -9'sd38;
	qsin_lut[3488] =  9'sd0;
	icos_lut[3488] = -9'sd37;
	qsin_lut[3489] = -9'sd7;
	icos_lut[3489] = -9'sd36;
	qsin_lut[3490] = -9'sd14;
	icos_lut[3490] = -9'sd34;
	qsin_lut[3491] = -9'sd21;
	icos_lut[3491] = -9'sd31;
	qsin_lut[3492] = -9'sd26;
	icos_lut[3492] = -9'sd26;
	qsin_lut[3493] = -9'sd31;
	icos_lut[3493] = -9'sd21;
	qsin_lut[3494] = -9'sd34;
	icos_lut[3494] = -9'sd14;
	qsin_lut[3495] = -9'sd36;
	icos_lut[3495] = -9'sd7;
	qsin_lut[3496] = -9'sd37;
	icos_lut[3496] = -9'sd0;
	qsin_lut[3497] = -9'sd36;
	icos_lut[3497] =  9'sd7;
	qsin_lut[3498] = -9'sd34;
	icos_lut[3498] =  9'sd14;
	qsin_lut[3499] = -9'sd31;
	icos_lut[3499] =  9'sd21;
	qsin_lut[3500] = -9'sd26;
	icos_lut[3500] =  9'sd26;
	qsin_lut[3501] = -9'sd21;
	icos_lut[3501] =  9'sd31;
	qsin_lut[3502] = -9'sd14;
	icos_lut[3502] =  9'sd34;
	qsin_lut[3503] = -9'sd7;
	icos_lut[3503] =  9'sd36;
	qsin_lut[3504] = -9'sd0;
	icos_lut[3504] =  9'sd37;
	qsin_lut[3505] =  9'sd7;
	icos_lut[3505] =  9'sd36;
	qsin_lut[3506] =  9'sd14;
	icos_lut[3506] =  9'sd34;
	qsin_lut[3507] =  9'sd21;
	icos_lut[3507] =  9'sd31;
	qsin_lut[3508] =  9'sd26;
	icos_lut[3508] =  9'sd26;
	qsin_lut[3509] =  9'sd31;
	icos_lut[3509] =  9'sd21;
	qsin_lut[3510] =  9'sd34;
	icos_lut[3510] =  9'sd14;
	qsin_lut[3511] =  9'sd36;
	icos_lut[3511] =  9'sd7;
	qsin_lut[3512] =  9'sd37;
	icos_lut[3512] =  9'sd0;
	qsin_lut[3513] =  9'sd36;
	icos_lut[3513] = -9'sd7;
	qsin_lut[3514] =  9'sd34;
	icos_lut[3514] = -9'sd14;
	qsin_lut[3515] =  9'sd31;
	icos_lut[3515] = -9'sd21;
	qsin_lut[3516] =  9'sd26;
	icos_lut[3516] = -9'sd26;
	qsin_lut[3517] =  9'sd21;
	icos_lut[3517] = -9'sd31;
	qsin_lut[3518] =  9'sd14;
	icos_lut[3518] = -9'sd34;
	qsin_lut[3519] =  9'sd7;
	icos_lut[3519] = -9'sd36;
	qsin_lut[3520] =  9'sd0;
	icos_lut[3520] = -9'sd35;
	qsin_lut[3521] = -9'sd7;
	icos_lut[3521] = -9'sd34;
	qsin_lut[3522] = -9'sd13;
	icos_lut[3522] = -9'sd32;
	qsin_lut[3523] = -9'sd19;
	icos_lut[3523] = -9'sd29;
	qsin_lut[3524] = -9'sd25;
	icos_lut[3524] = -9'sd25;
	qsin_lut[3525] = -9'sd29;
	icos_lut[3525] = -9'sd19;
	qsin_lut[3526] = -9'sd32;
	icos_lut[3526] = -9'sd13;
	qsin_lut[3527] = -9'sd34;
	icos_lut[3527] = -9'sd7;
	qsin_lut[3528] = -9'sd35;
	icos_lut[3528] = -9'sd0;
	qsin_lut[3529] = -9'sd34;
	icos_lut[3529] =  9'sd7;
	qsin_lut[3530] = -9'sd32;
	icos_lut[3530] =  9'sd13;
	qsin_lut[3531] = -9'sd29;
	icos_lut[3531] =  9'sd19;
	qsin_lut[3532] = -9'sd25;
	icos_lut[3532] =  9'sd25;
	qsin_lut[3533] = -9'sd19;
	icos_lut[3533] =  9'sd29;
	qsin_lut[3534] = -9'sd13;
	icos_lut[3534] =  9'sd32;
	qsin_lut[3535] = -9'sd7;
	icos_lut[3535] =  9'sd34;
	qsin_lut[3536] = -9'sd0;
	icos_lut[3536] =  9'sd35;
	qsin_lut[3537] =  9'sd7;
	icos_lut[3537] =  9'sd34;
	qsin_lut[3538] =  9'sd13;
	icos_lut[3538] =  9'sd32;
	qsin_lut[3539] =  9'sd19;
	icos_lut[3539] =  9'sd29;
	qsin_lut[3540] =  9'sd25;
	icos_lut[3540] =  9'sd25;
	qsin_lut[3541] =  9'sd29;
	icos_lut[3541] =  9'sd19;
	qsin_lut[3542] =  9'sd32;
	icos_lut[3542] =  9'sd13;
	qsin_lut[3543] =  9'sd34;
	icos_lut[3543] =  9'sd7;
	qsin_lut[3544] =  9'sd35;
	icos_lut[3544] =  9'sd0;
	qsin_lut[3545] =  9'sd34;
	icos_lut[3545] = -9'sd7;
	qsin_lut[3546] =  9'sd32;
	icos_lut[3546] = -9'sd13;
	qsin_lut[3547] =  9'sd29;
	icos_lut[3547] = -9'sd19;
	qsin_lut[3548] =  9'sd25;
	icos_lut[3548] = -9'sd25;
	qsin_lut[3549] =  9'sd19;
	icos_lut[3549] = -9'sd29;
	qsin_lut[3550] =  9'sd13;
	icos_lut[3550] = -9'sd32;
	qsin_lut[3551] =  9'sd7;
	icos_lut[3551] = -9'sd34;
	qsin_lut[3552] =  9'sd0;
	icos_lut[3552] = -9'sd33;
	qsin_lut[3553] = -9'sd6;
	icos_lut[3553] = -9'sd32;
	qsin_lut[3554] = -9'sd13;
	icos_lut[3554] = -9'sd30;
	qsin_lut[3555] = -9'sd18;
	icos_lut[3555] = -9'sd27;
	qsin_lut[3556] = -9'sd23;
	icos_lut[3556] = -9'sd23;
	qsin_lut[3557] = -9'sd27;
	icos_lut[3557] = -9'sd18;
	qsin_lut[3558] = -9'sd30;
	icos_lut[3558] = -9'sd13;
	qsin_lut[3559] = -9'sd32;
	icos_lut[3559] = -9'sd6;
	qsin_lut[3560] = -9'sd33;
	icos_lut[3560] = -9'sd0;
	qsin_lut[3561] = -9'sd32;
	icos_lut[3561] =  9'sd6;
	qsin_lut[3562] = -9'sd30;
	icos_lut[3562] =  9'sd13;
	qsin_lut[3563] = -9'sd27;
	icos_lut[3563] =  9'sd18;
	qsin_lut[3564] = -9'sd23;
	icos_lut[3564] =  9'sd23;
	qsin_lut[3565] = -9'sd18;
	icos_lut[3565] =  9'sd27;
	qsin_lut[3566] = -9'sd13;
	icos_lut[3566] =  9'sd30;
	qsin_lut[3567] = -9'sd6;
	icos_lut[3567] =  9'sd32;
	qsin_lut[3568] = -9'sd0;
	icos_lut[3568] =  9'sd33;
	qsin_lut[3569] =  9'sd6;
	icos_lut[3569] =  9'sd32;
	qsin_lut[3570] =  9'sd13;
	icos_lut[3570] =  9'sd30;
	qsin_lut[3571] =  9'sd18;
	icos_lut[3571] =  9'sd27;
	qsin_lut[3572] =  9'sd23;
	icos_lut[3572] =  9'sd23;
	qsin_lut[3573] =  9'sd27;
	icos_lut[3573] =  9'sd18;
	qsin_lut[3574] =  9'sd30;
	icos_lut[3574] =  9'sd13;
	qsin_lut[3575] =  9'sd32;
	icos_lut[3575] =  9'sd6;
	qsin_lut[3576] =  9'sd33;
	icos_lut[3576] =  9'sd0;
	qsin_lut[3577] =  9'sd32;
	icos_lut[3577] = -9'sd6;
	qsin_lut[3578] =  9'sd30;
	icos_lut[3578] = -9'sd13;
	qsin_lut[3579] =  9'sd27;
	icos_lut[3579] = -9'sd18;
	qsin_lut[3580] =  9'sd23;
	icos_lut[3580] = -9'sd23;
	qsin_lut[3581] =  9'sd18;
	icos_lut[3581] = -9'sd27;
	qsin_lut[3582] =  9'sd13;
	icos_lut[3582] = -9'sd30;
	qsin_lut[3583] =  9'sd6;
	icos_lut[3583] = -9'sd32;
	qsin_lut[3584] =  9'sd0;
	icos_lut[3584] = -9'sd31;
	qsin_lut[3585] = -9'sd6;
	icos_lut[3585] = -9'sd30;
	qsin_lut[3586] = -9'sd12;
	icos_lut[3586] = -9'sd29;
	qsin_lut[3587] = -9'sd17;
	icos_lut[3587] = -9'sd26;
	qsin_lut[3588] = -9'sd22;
	icos_lut[3588] = -9'sd22;
	qsin_lut[3589] = -9'sd26;
	icos_lut[3589] = -9'sd17;
	qsin_lut[3590] = -9'sd29;
	icos_lut[3590] = -9'sd12;
	qsin_lut[3591] = -9'sd30;
	icos_lut[3591] = -9'sd6;
	qsin_lut[3592] = -9'sd31;
	icos_lut[3592] = -9'sd0;
	qsin_lut[3593] = -9'sd30;
	icos_lut[3593] =  9'sd6;
	qsin_lut[3594] = -9'sd29;
	icos_lut[3594] =  9'sd12;
	qsin_lut[3595] = -9'sd26;
	icos_lut[3595] =  9'sd17;
	qsin_lut[3596] = -9'sd22;
	icos_lut[3596] =  9'sd22;
	qsin_lut[3597] = -9'sd17;
	icos_lut[3597] =  9'sd26;
	qsin_lut[3598] = -9'sd12;
	icos_lut[3598] =  9'sd29;
	qsin_lut[3599] = -9'sd6;
	icos_lut[3599] =  9'sd30;
	qsin_lut[3600] = -9'sd0;
	icos_lut[3600] =  9'sd31;
	qsin_lut[3601] =  9'sd6;
	icos_lut[3601] =  9'sd30;
	qsin_lut[3602] =  9'sd12;
	icos_lut[3602] =  9'sd29;
	qsin_lut[3603] =  9'sd17;
	icos_lut[3603] =  9'sd26;
	qsin_lut[3604] =  9'sd22;
	icos_lut[3604] =  9'sd22;
	qsin_lut[3605] =  9'sd26;
	icos_lut[3605] =  9'sd17;
	qsin_lut[3606] =  9'sd29;
	icos_lut[3606] =  9'sd12;
	qsin_lut[3607] =  9'sd30;
	icos_lut[3607] =  9'sd6;
	qsin_lut[3608] =  9'sd31;
	icos_lut[3608] =  9'sd0;
	qsin_lut[3609] =  9'sd30;
	icos_lut[3609] = -9'sd6;
	qsin_lut[3610] =  9'sd29;
	icos_lut[3610] = -9'sd12;
	qsin_lut[3611] =  9'sd26;
	icos_lut[3611] = -9'sd17;
	qsin_lut[3612] =  9'sd22;
	icos_lut[3612] = -9'sd22;
	qsin_lut[3613] =  9'sd17;
	icos_lut[3613] = -9'sd26;
	qsin_lut[3614] =  9'sd12;
	icos_lut[3614] = -9'sd29;
	qsin_lut[3615] =  9'sd6;
	icos_lut[3615] = -9'sd30;
	qsin_lut[3616] =  9'sd0;
	icos_lut[3616] = -9'sd29;
	qsin_lut[3617] = -9'sd6;
	icos_lut[3617] = -9'sd28;
	qsin_lut[3618] = -9'sd11;
	icos_lut[3618] = -9'sd27;
	qsin_lut[3619] = -9'sd16;
	icos_lut[3619] = -9'sd24;
	qsin_lut[3620] = -9'sd21;
	icos_lut[3620] = -9'sd21;
	qsin_lut[3621] = -9'sd24;
	icos_lut[3621] = -9'sd16;
	qsin_lut[3622] = -9'sd27;
	icos_lut[3622] = -9'sd11;
	qsin_lut[3623] = -9'sd28;
	icos_lut[3623] = -9'sd6;
	qsin_lut[3624] = -9'sd29;
	icos_lut[3624] = -9'sd0;
	qsin_lut[3625] = -9'sd28;
	icos_lut[3625] =  9'sd6;
	qsin_lut[3626] = -9'sd27;
	icos_lut[3626] =  9'sd11;
	qsin_lut[3627] = -9'sd24;
	icos_lut[3627] =  9'sd16;
	qsin_lut[3628] = -9'sd21;
	icos_lut[3628] =  9'sd21;
	qsin_lut[3629] = -9'sd16;
	icos_lut[3629] =  9'sd24;
	qsin_lut[3630] = -9'sd11;
	icos_lut[3630] =  9'sd27;
	qsin_lut[3631] = -9'sd6;
	icos_lut[3631] =  9'sd28;
	qsin_lut[3632] = -9'sd0;
	icos_lut[3632] =  9'sd29;
	qsin_lut[3633] =  9'sd6;
	icos_lut[3633] =  9'sd28;
	qsin_lut[3634] =  9'sd11;
	icos_lut[3634] =  9'sd27;
	qsin_lut[3635] =  9'sd16;
	icos_lut[3635] =  9'sd24;
	qsin_lut[3636] =  9'sd21;
	icos_lut[3636] =  9'sd21;
	qsin_lut[3637] =  9'sd24;
	icos_lut[3637] =  9'sd16;
	qsin_lut[3638] =  9'sd27;
	icos_lut[3638] =  9'sd11;
	qsin_lut[3639] =  9'sd28;
	icos_lut[3639] =  9'sd6;
	qsin_lut[3640] =  9'sd29;
	icos_lut[3640] =  9'sd0;
	qsin_lut[3641] =  9'sd28;
	icos_lut[3641] = -9'sd6;
	qsin_lut[3642] =  9'sd27;
	icos_lut[3642] = -9'sd11;
	qsin_lut[3643] =  9'sd24;
	icos_lut[3643] = -9'sd16;
	qsin_lut[3644] =  9'sd21;
	icos_lut[3644] = -9'sd21;
	qsin_lut[3645] =  9'sd16;
	icos_lut[3645] = -9'sd24;
	qsin_lut[3646] =  9'sd11;
	icos_lut[3646] = -9'sd27;
	qsin_lut[3647] =  9'sd6;
	icos_lut[3647] = -9'sd28;
	qsin_lut[3648] =  9'sd0;
	icos_lut[3648] = -9'sd27;
	qsin_lut[3649] = -9'sd5;
	icos_lut[3649] = -9'sd26;
	qsin_lut[3650] = -9'sd10;
	icos_lut[3650] = -9'sd25;
	qsin_lut[3651] = -9'sd15;
	icos_lut[3651] = -9'sd22;
	qsin_lut[3652] = -9'sd19;
	icos_lut[3652] = -9'sd19;
	qsin_lut[3653] = -9'sd22;
	icos_lut[3653] = -9'sd15;
	qsin_lut[3654] = -9'sd25;
	icos_lut[3654] = -9'sd10;
	qsin_lut[3655] = -9'sd26;
	icos_lut[3655] = -9'sd5;
	qsin_lut[3656] = -9'sd27;
	icos_lut[3656] = -9'sd0;
	qsin_lut[3657] = -9'sd26;
	icos_lut[3657] =  9'sd5;
	qsin_lut[3658] = -9'sd25;
	icos_lut[3658] =  9'sd10;
	qsin_lut[3659] = -9'sd22;
	icos_lut[3659] =  9'sd15;
	qsin_lut[3660] = -9'sd19;
	icos_lut[3660] =  9'sd19;
	qsin_lut[3661] = -9'sd15;
	icos_lut[3661] =  9'sd22;
	qsin_lut[3662] = -9'sd10;
	icos_lut[3662] =  9'sd25;
	qsin_lut[3663] = -9'sd5;
	icos_lut[3663] =  9'sd26;
	qsin_lut[3664] = -9'sd0;
	icos_lut[3664] =  9'sd27;
	qsin_lut[3665] =  9'sd5;
	icos_lut[3665] =  9'sd26;
	qsin_lut[3666] =  9'sd10;
	icos_lut[3666] =  9'sd25;
	qsin_lut[3667] =  9'sd15;
	icos_lut[3667] =  9'sd22;
	qsin_lut[3668] =  9'sd19;
	icos_lut[3668] =  9'sd19;
	qsin_lut[3669] =  9'sd22;
	icos_lut[3669] =  9'sd15;
	qsin_lut[3670] =  9'sd25;
	icos_lut[3670] =  9'sd10;
	qsin_lut[3671] =  9'sd26;
	icos_lut[3671] =  9'sd5;
	qsin_lut[3672] =  9'sd27;
	icos_lut[3672] =  9'sd0;
	qsin_lut[3673] =  9'sd26;
	icos_lut[3673] = -9'sd5;
	qsin_lut[3674] =  9'sd25;
	icos_lut[3674] = -9'sd10;
	qsin_lut[3675] =  9'sd22;
	icos_lut[3675] = -9'sd15;
	qsin_lut[3676] =  9'sd19;
	icos_lut[3676] = -9'sd19;
	qsin_lut[3677] =  9'sd15;
	icos_lut[3677] = -9'sd22;
	qsin_lut[3678] =  9'sd10;
	icos_lut[3678] = -9'sd25;
	qsin_lut[3679] =  9'sd5;
	icos_lut[3679] = -9'sd26;
	qsin_lut[3680] =  9'sd0;
	icos_lut[3680] = -9'sd25;
	qsin_lut[3681] = -9'sd5;
	icos_lut[3681] = -9'sd25;
	qsin_lut[3682] = -9'sd10;
	icos_lut[3682] = -9'sd23;
	qsin_lut[3683] = -9'sd14;
	icos_lut[3683] = -9'sd21;
	qsin_lut[3684] = -9'sd18;
	icos_lut[3684] = -9'sd18;
	qsin_lut[3685] = -9'sd21;
	icos_lut[3685] = -9'sd14;
	qsin_lut[3686] = -9'sd23;
	icos_lut[3686] = -9'sd10;
	qsin_lut[3687] = -9'sd25;
	icos_lut[3687] = -9'sd5;
	qsin_lut[3688] = -9'sd25;
	icos_lut[3688] = -9'sd0;
	qsin_lut[3689] = -9'sd25;
	icos_lut[3689] =  9'sd5;
	qsin_lut[3690] = -9'sd23;
	icos_lut[3690] =  9'sd10;
	qsin_lut[3691] = -9'sd21;
	icos_lut[3691] =  9'sd14;
	qsin_lut[3692] = -9'sd18;
	icos_lut[3692] =  9'sd18;
	qsin_lut[3693] = -9'sd14;
	icos_lut[3693] =  9'sd21;
	qsin_lut[3694] = -9'sd10;
	icos_lut[3694] =  9'sd23;
	qsin_lut[3695] = -9'sd5;
	icos_lut[3695] =  9'sd25;
	qsin_lut[3696] = -9'sd0;
	icos_lut[3696] =  9'sd25;
	qsin_lut[3697] =  9'sd5;
	icos_lut[3697] =  9'sd25;
	qsin_lut[3698] =  9'sd10;
	icos_lut[3698] =  9'sd23;
	qsin_lut[3699] =  9'sd14;
	icos_lut[3699] =  9'sd21;
	qsin_lut[3700] =  9'sd18;
	icos_lut[3700] =  9'sd18;
	qsin_lut[3701] =  9'sd21;
	icos_lut[3701] =  9'sd14;
	qsin_lut[3702] =  9'sd23;
	icos_lut[3702] =  9'sd10;
	qsin_lut[3703] =  9'sd25;
	icos_lut[3703] =  9'sd5;
	qsin_lut[3704] =  9'sd25;
	icos_lut[3704] =  9'sd0;
	qsin_lut[3705] =  9'sd25;
	icos_lut[3705] = -9'sd5;
	qsin_lut[3706] =  9'sd23;
	icos_lut[3706] = -9'sd10;
	qsin_lut[3707] =  9'sd21;
	icos_lut[3707] = -9'sd14;
	qsin_lut[3708] =  9'sd18;
	icos_lut[3708] = -9'sd18;
	qsin_lut[3709] =  9'sd14;
	icos_lut[3709] = -9'sd21;
	qsin_lut[3710] =  9'sd10;
	icos_lut[3710] = -9'sd23;
	qsin_lut[3711] =  9'sd5;
	icos_lut[3711] = -9'sd25;
	qsin_lut[3712] =  9'sd0;
	icos_lut[3712] = -9'sd23;
	qsin_lut[3713] = -9'sd4;
	icos_lut[3713] = -9'sd23;
	qsin_lut[3714] = -9'sd9;
	icos_lut[3714] = -9'sd21;
	qsin_lut[3715] = -9'sd13;
	icos_lut[3715] = -9'sd19;
	qsin_lut[3716] = -9'sd16;
	icos_lut[3716] = -9'sd16;
	qsin_lut[3717] = -9'sd19;
	icos_lut[3717] = -9'sd13;
	qsin_lut[3718] = -9'sd21;
	icos_lut[3718] = -9'sd9;
	qsin_lut[3719] = -9'sd23;
	icos_lut[3719] = -9'sd4;
	qsin_lut[3720] = -9'sd23;
	icos_lut[3720] = -9'sd0;
	qsin_lut[3721] = -9'sd23;
	icos_lut[3721] =  9'sd4;
	qsin_lut[3722] = -9'sd21;
	icos_lut[3722] =  9'sd9;
	qsin_lut[3723] = -9'sd19;
	icos_lut[3723] =  9'sd13;
	qsin_lut[3724] = -9'sd16;
	icos_lut[3724] =  9'sd16;
	qsin_lut[3725] = -9'sd13;
	icos_lut[3725] =  9'sd19;
	qsin_lut[3726] = -9'sd9;
	icos_lut[3726] =  9'sd21;
	qsin_lut[3727] = -9'sd4;
	icos_lut[3727] =  9'sd23;
	qsin_lut[3728] = -9'sd0;
	icos_lut[3728] =  9'sd23;
	qsin_lut[3729] =  9'sd4;
	icos_lut[3729] =  9'sd23;
	qsin_lut[3730] =  9'sd9;
	icos_lut[3730] =  9'sd21;
	qsin_lut[3731] =  9'sd13;
	icos_lut[3731] =  9'sd19;
	qsin_lut[3732] =  9'sd16;
	icos_lut[3732] =  9'sd16;
	qsin_lut[3733] =  9'sd19;
	icos_lut[3733] =  9'sd13;
	qsin_lut[3734] =  9'sd21;
	icos_lut[3734] =  9'sd9;
	qsin_lut[3735] =  9'sd23;
	icos_lut[3735] =  9'sd4;
	qsin_lut[3736] =  9'sd23;
	icos_lut[3736] =  9'sd0;
	qsin_lut[3737] =  9'sd23;
	icos_lut[3737] = -9'sd4;
	qsin_lut[3738] =  9'sd21;
	icos_lut[3738] = -9'sd9;
	qsin_lut[3739] =  9'sd19;
	icos_lut[3739] = -9'sd13;
	qsin_lut[3740] =  9'sd16;
	icos_lut[3740] = -9'sd16;
	qsin_lut[3741] =  9'sd13;
	icos_lut[3741] = -9'sd19;
	qsin_lut[3742] =  9'sd9;
	icos_lut[3742] = -9'sd21;
	qsin_lut[3743] =  9'sd4;
	icos_lut[3743] = -9'sd23;
	qsin_lut[3744] =  9'sd0;
	icos_lut[3744] = -9'sd21;
	qsin_lut[3745] = -9'sd4;
	icos_lut[3745] = -9'sd21;
	qsin_lut[3746] = -9'sd8;
	icos_lut[3746] = -9'sd19;
	qsin_lut[3747] = -9'sd12;
	icos_lut[3747] = -9'sd17;
	qsin_lut[3748] = -9'sd15;
	icos_lut[3748] = -9'sd15;
	qsin_lut[3749] = -9'sd17;
	icos_lut[3749] = -9'sd12;
	qsin_lut[3750] = -9'sd19;
	icos_lut[3750] = -9'sd8;
	qsin_lut[3751] = -9'sd21;
	icos_lut[3751] = -9'sd4;
	qsin_lut[3752] = -9'sd21;
	icos_lut[3752] = -9'sd0;
	qsin_lut[3753] = -9'sd21;
	icos_lut[3753] =  9'sd4;
	qsin_lut[3754] = -9'sd19;
	icos_lut[3754] =  9'sd8;
	qsin_lut[3755] = -9'sd17;
	icos_lut[3755] =  9'sd12;
	qsin_lut[3756] = -9'sd15;
	icos_lut[3756] =  9'sd15;
	qsin_lut[3757] = -9'sd12;
	icos_lut[3757] =  9'sd17;
	qsin_lut[3758] = -9'sd8;
	icos_lut[3758] =  9'sd19;
	qsin_lut[3759] = -9'sd4;
	icos_lut[3759] =  9'sd21;
	qsin_lut[3760] = -9'sd0;
	icos_lut[3760] =  9'sd21;
	qsin_lut[3761] =  9'sd4;
	icos_lut[3761] =  9'sd21;
	qsin_lut[3762] =  9'sd8;
	icos_lut[3762] =  9'sd19;
	qsin_lut[3763] =  9'sd12;
	icos_lut[3763] =  9'sd17;
	qsin_lut[3764] =  9'sd15;
	icos_lut[3764] =  9'sd15;
	qsin_lut[3765] =  9'sd17;
	icos_lut[3765] =  9'sd12;
	qsin_lut[3766] =  9'sd19;
	icos_lut[3766] =  9'sd8;
	qsin_lut[3767] =  9'sd21;
	icos_lut[3767] =  9'sd4;
	qsin_lut[3768] =  9'sd21;
	icos_lut[3768] =  9'sd0;
	qsin_lut[3769] =  9'sd21;
	icos_lut[3769] = -9'sd4;
	qsin_lut[3770] =  9'sd19;
	icos_lut[3770] = -9'sd8;
	qsin_lut[3771] =  9'sd17;
	icos_lut[3771] = -9'sd12;
	qsin_lut[3772] =  9'sd15;
	icos_lut[3772] = -9'sd15;
	qsin_lut[3773] =  9'sd12;
	icos_lut[3773] = -9'sd17;
	qsin_lut[3774] =  9'sd8;
	icos_lut[3774] = -9'sd19;
	qsin_lut[3775] =  9'sd4;
	icos_lut[3775] = -9'sd21;
	qsin_lut[3776] =  9'sd0;
	icos_lut[3776] = -9'sd19;
	qsin_lut[3777] = -9'sd4;
	icos_lut[3777] = -9'sd19;
	qsin_lut[3778] = -9'sd7;
	icos_lut[3778] = -9'sd18;
	qsin_lut[3779] = -9'sd11;
	icos_lut[3779] = -9'sd16;
	qsin_lut[3780] = -9'sd13;
	icos_lut[3780] = -9'sd13;
	qsin_lut[3781] = -9'sd16;
	icos_lut[3781] = -9'sd11;
	qsin_lut[3782] = -9'sd18;
	icos_lut[3782] = -9'sd7;
	qsin_lut[3783] = -9'sd19;
	icos_lut[3783] = -9'sd4;
	qsin_lut[3784] = -9'sd19;
	icos_lut[3784] = -9'sd0;
	qsin_lut[3785] = -9'sd19;
	icos_lut[3785] =  9'sd4;
	qsin_lut[3786] = -9'sd18;
	icos_lut[3786] =  9'sd7;
	qsin_lut[3787] = -9'sd16;
	icos_lut[3787] =  9'sd11;
	qsin_lut[3788] = -9'sd13;
	icos_lut[3788] =  9'sd13;
	qsin_lut[3789] = -9'sd11;
	icos_lut[3789] =  9'sd16;
	qsin_lut[3790] = -9'sd7;
	icos_lut[3790] =  9'sd18;
	qsin_lut[3791] = -9'sd4;
	icos_lut[3791] =  9'sd19;
	qsin_lut[3792] = -9'sd0;
	icos_lut[3792] =  9'sd19;
	qsin_lut[3793] =  9'sd4;
	icos_lut[3793] =  9'sd19;
	qsin_lut[3794] =  9'sd7;
	icos_lut[3794] =  9'sd18;
	qsin_lut[3795] =  9'sd11;
	icos_lut[3795] =  9'sd16;
	qsin_lut[3796] =  9'sd13;
	icos_lut[3796] =  9'sd13;
	qsin_lut[3797] =  9'sd16;
	icos_lut[3797] =  9'sd11;
	qsin_lut[3798] =  9'sd18;
	icos_lut[3798] =  9'sd7;
	qsin_lut[3799] =  9'sd19;
	icos_lut[3799] =  9'sd4;
	qsin_lut[3800] =  9'sd19;
	icos_lut[3800] =  9'sd0;
	qsin_lut[3801] =  9'sd19;
	icos_lut[3801] = -9'sd4;
	qsin_lut[3802] =  9'sd18;
	icos_lut[3802] = -9'sd7;
	qsin_lut[3803] =  9'sd16;
	icos_lut[3803] = -9'sd11;
	qsin_lut[3804] =  9'sd13;
	icos_lut[3804] = -9'sd13;
	qsin_lut[3805] =  9'sd11;
	icos_lut[3805] = -9'sd16;
	qsin_lut[3806] =  9'sd7;
	icos_lut[3806] = -9'sd18;
	qsin_lut[3807] =  9'sd4;
	icos_lut[3807] = -9'sd19;
	qsin_lut[3808] =  9'sd0;
	icos_lut[3808] = -9'sd17;
	qsin_lut[3809] = -9'sd3;
	icos_lut[3809] = -9'sd17;
	qsin_lut[3810] = -9'sd7;
	icos_lut[3810] = -9'sd16;
	qsin_lut[3811] = -9'sd9;
	icos_lut[3811] = -9'sd14;
	qsin_lut[3812] = -9'sd12;
	icos_lut[3812] = -9'sd12;
	qsin_lut[3813] = -9'sd14;
	icos_lut[3813] = -9'sd9;
	qsin_lut[3814] = -9'sd16;
	icos_lut[3814] = -9'sd7;
	qsin_lut[3815] = -9'sd17;
	icos_lut[3815] = -9'sd3;
	qsin_lut[3816] = -9'sd17;
	icos_lut[3816] = -9'sd0;
	qsin_lut[3817] = -9'sd17;
	icos_lut[3817] =  9'sd3;
	qsin_lut[3818] = -9'sd16;
	icos_lut[3818] =  9'sd7;
	qsin_lut[3819] = -9'sd14;
	icos_lut[3819] =  9'sd9;
	qsin_lut[3820] = -9'sd12;
	icos_lut[3820] =  9'sd12;
	qsin_lut[3821] = -9'sd9;
	icos_lut[3821] =  9'sd14;
	qsin_lut[3822] = -9'sd7;
	icos_lut[3822] =  9'sd16;
	qsin_lut[3823] = -9'sd3;
	icos_lut[3823] =  9'sd17;
	qsin_lut[3824] = -9'sd0;
	icos_lut[3824] =  9'sd17;
	qsin_lut[3825] =  9'sd3;
	icos_lut[3825] =  9'sd17;
	qsin_lut[3826] =  9'sd7;
	icos_lut[3826] =  9'sd16;
	qsin_lut[3827] =  9'sd9;
	icos_lut[3827] =  9'sd14;
	qsin_lut[3828] =  9'sd12;
	icos_lut[3828] =  9'sd12;
	qsin_lut[3829] =  9'sd14;
	icos_lut[3829] =  9'sd9;
	qsin_lut[3830] =  9'sd16;
	icos_lut[3830] =  9'sd7;
	qsin_lut[3831] =  9'sd17;
	icos_lut[3831] =  9'sd3;
	qsin_lut[3832] =  9'sd17;
	icos_lut[3832] =  9'sd0;
	qsin_lut[3833] =  9'sd17;
	icos_lut[3833] = -9'sd3;
	qsin_lut[3834] =  9'sd16;
	icos_lut[3834] = -9'sd7;
	qsin_lut[3835] =  9'sd14;
	icos_lut[3835] = -9'sd9;
	qsin_lut[3836] =  9'sd12;
	icos_lut[3836] = -9'sd12;
	qsin_lut[3837] =  9'sd9;
	icos_lut[3837] = -9'sd14;
	qsin_lut[3838] =  9'sd7;
	icos_lut[3838] = -9'sd16;
	qsin_lut[3839] =  9'sd3;
	icos_lut[3839] = -9'sd17;
	qsin_lut[3840] =  9'sd0;
	icos_lut[3840] = -9'sd15;
	qsin_lut[3841] = -9'sd3;
	icos_lut[3841] = -9'sd15;
	qsin_lut[3842] = -9'sd6;
	icos_lut[3842] = -9'sd14;
	qsin_lut[3843] = -9'sd8;
	icos_lut[3843] = -9'sd12;
	qsin_lut[3844] = -9'sd11;
	icos_lut[3844] = -9'sd11;
	qsin_lut[3845] = -9'sd12;
	icos_lut[3845] = -9'sd8;
	qsin_lut[3846] = -9'sd14;
	icos_lut[3846] = -9'sd6;
	qsin_lut[3847] = -9'sd15;
	icos_lut[3847] = -9'sd3;
	qsin_lut[3848] = -9'sd15;
	icos_lut[3848] = -9'sd0;
	qsin_lut[3849] = -9'sd15;
	icos_lut[3849] =  9'sd3;
	qsin_lut[3850] = -9'sd14;
	icos_lut[3850] =  9'sd6;
	qsin_lut[3851] = -9'sd12;
	icos_lut[3851] =  9'sd8;
	qsin_lut[3852] = -9'sd11;
	icos_lut[3852] =  9'sd11;
	qsin_lut[3853] = -9'sd8;
	icos_lut[3853] =  9'sd12;
	qsin_lut[3854] = -9'sd6;
	icos_lut[3854] =  9'sd14;
	qsin_lut[3855] = -9'sd3;
	icos_lut[3855] =  9'sd15;
	qsin_lut[3856] = -9'sd0;
	icos_lut[3856] =  9'sd15;
	qsin_lut[3857] =  9'sd3;
	icos_lut[3857] =  9'sd15;
	qsin_lut[3858] =  9'sd6;
	icos_lut[3858] =  9'sd14;
	qsin_lut[3859] =  9'sd8;
	icos_lut[3859] =  9'sd12;
	qsin_lut[3860] =  9'sd11;
	icos_lut[3860] =  9'sd11;
	qsin_lut[3861] =  9'sd12;
	icos_lut[3861] =  9'sd8;
	qsin_lut[3862] =  9'sd14;
	icos_lut[3862] =  9'sd6;
	qsin_lut[3863] =  9'sd15;
	icos_lut[3863] =  9'sd3;
	qsin_lut[3864] =  9'sd15;
	icos_lut[3864] =  9'sd0;
	qsin_lut[3865] =  9'sd15;
	icos_lut[3865] = -9'sd3;
	qsin_lut[3866] =  9'sd14;
	icos_lut[3866] = -9'sd6;
	qsin_lut[3867] =  9'sd12;
	icos_lut[3867] = -9'sd8;
	qsin_lut[3868] =  9'sd11;
	icos_lut[3868] = -9'sd11;
	qsin_lut[3869] =  9'sd8;
	icos_lut[3869] = -9'sd12;
	qsin_lut[3870] =  9'sd6;
	icos_lut[3870] = -9'sd14;
	qsin_lut[3871] =  9'sd3;
	icos_lut[3871] = -9'sd15;
	qsin_lut[3872] =  9'sd0;
	icos_lut[3872] = -9'sd13;
	qsin_lut[3873] = -9'sd3;
	icos_lut[3873] = -9'sd13;
	qsin_lut[3874] = -9'sd5;
	icos_lut[3874] = -9'sd12;
	qsin_lut[3875] = -9'sd7;
	icos_lut[3875] = -9'sd11;
	qsin_lut[3876] = -9'sd9;
	icos_lut[3876] = -9'sd9;
	qsin_lut[3877] = -9'sd11;
	icos_lut[3877] = -9'sd7;
	qsin_lut[3878] = -9'sd12;
	icos_lut[3878] = -9'sd5;
	qsin_lut[3879] = -9'sd13;
	icos_lut[3879] = -9'sd3;
	qsin_lut[3880] = -9'sd13;
	icos_lut[3880] = -9'sd0;
	qsin_lut[3881] = -9'sd13;
	icos_lut[3881] =  9'sd3;
	qsin_lut[3882] = -9'sd12;
	icos_lut[3882] =  9'sd5;
	qsin_lut[3883] = -9'sd11;
	icos_lut[3883] =  9'sd7;
	qsin_lut[3884] = -9'sd9;
	icos_lut[3884] =  9'sd9;
	qsin_lut[3885] = -9'sd7;
	icos_lut[3885] =  9'sd11;
	qsin_lut[3886] = -9'sd5;
	icos_lut[3886] =  9'sd12;
	qsin_lut[3887] = -9'sd3;
	icos_lut[3887] =  9'sd13;
	qsin_lut[3888] = -9'sd0;
	icos_lut[3888] =  9'sd13;
	qsin_lut[3889] =  9'sd3;
	icos_lut[3889] =  9'sd13;
	qsin_lut[3890] =  9'sd5;
	icos_lut[3890] =  9'sd12;
	qsin_lut[3891] =  9'sd7;
	icos_lut[3891] =  9'sd11;
	qsin_lut[3892] =  9'sd9;
	icos_lut[3892] =  9'sd9;
	qsin_lut[3893] =  9'sd11;
	icos_lut[3893] =  9'sd7;
	qsin_lut[3894] =  9'sd12;
	icos_lut[3894] =  9'sd5;
	qsin_lut[3895] =  9'sd13;
	icos_lut[3895] =  9'sd3;
	qsin_lut[3896] =  9'sd13;
	icos_lut[3896] =  9'sd0;
	qsin_lut[3897] =  9'sd13;
	icos_lut[3897] = -9'sd3;
	qsin_lut[3898] =  9'sd12;
	icos_lut[3898] = -9'sd5;
	qsin_lut[3899] =  9'sd11;
	icos_lut[3899] = -9'sd7;
	qsin_lut[3900] =  9'sd9;
	icos_lut[3900] = -9'sd9;
	qsin_lut[3901] =  9'sd7;
	icos_lut[3901] = -9'sd11;
	qsin_lut[3902] =  9'sd5;
	icos_lut[3902] = -9'sd12;
	qsin_lut[3903] =  9'sd3;
	icos_lut[3903] = -9'sd13;
	qsin_lut[3904] =  9'sd0;
	icos_lut[3904] = -9'sd11;
	qsin_lut[3905] = -9'sd2;
	icos_lut[3905] = -9'sd11;
	qsin_lut[3906] = -9'sd4;
	icos_lut[3906] = -9'sd10;
	qsin_lut[3907] = -9'sd6;
	icos_lut[3907] = -9'sd9;
	qsin_lut[3908] = -9'sd8;
	icos_lut[3908] = -9'sd8;
	qsin_lut[3909] = -9'sd9;
	icos_lut[3909] = -9'sd6;
	qsin_lut[3910] = -9'sd10;
	icos_lut[3910] = -9'sd4;
	qsin_lut[3911] = -9'sd11;
	icos_lut[3911] = -9'sd2;
	qsin_lut[3912] = -9'sd11;
	icos_lut[3912] = -9'sd0;
	qsin_lut[3913] = -9'sd11;
	icos_lut[3913] =  9'sd2;
	qsin_lut[3914] = -9'sd10;
	icos_lut[3914] =  9'sd4;
	qsin_lut[3915] = -9'sd9;
	icos_lut[3915] =  9'sd6;
	qsin_lut[3916] = -9'sd8;
	icos_lut[3916] =  9'sd8;
	qsin_lut[3917] = -9'sd6;
	icos_lut[3917] =  9'sd9;
	qsin_lut[3918] = -9'sd4;
	icos_lut[3918] =  9'sd10;
	qsin_lut[3919] = -9'sd2;
	icos_lut[3919] =  9'sd11;
	qsin_lut[3920] = -9'sd0;
	icos_lut[3920] =  9'sd11;
	qsin_lut[3921] =  9'sd2;
	icos_lut[3921] =  9'sd11;
	qsin_lut[3922] =  9'sd4;
	icos_lut[3922] =  9'sd10;
	qsin_lut[3923] =  9'sd6;
	icos_lut[3923] =  9'sd9;
	qsin_lut[3924] =  9'sd8;
	icos_lut[3924] =  9'sd8;
	qsin_lut[3925] =  9'sd9;
	icos_lut[3925] =  9'sd6;
	qsin_lut[3926] =  9'sd10;
	icos_lut[3926] =  9'sd4;
	qsin_lut[3927] =  9'sd11;
	icos_lut[3927] =  9'sd2;
	qsin_lut[3928] =  9'sd11;
	icos_lut[3928] =  9'sd0;
	qsin_lut[3929] =  9'sd11;
	icos_lut[3929] = -9'sd2;
	qsin_lut[3930] =  9'sd10;
	icos_lut[3930] = -9'sd4;
	qsin_lut[3931] =  9'sd9;
	icos_lut[3931] = -9'sd6;
	qsin_lut[3932] =  9'sd8;
	icos_lut[3932] = -9'sd8;
	qsin_lut[3933] =  9'sd6;
	icos_lut[3933] = -9'sd9;
	qsin_lut[3934] =  9'sd4;
	icos_lut[3934] = -9'sd10;
	qsin_lut[3935] =  9'sd2;
	icos_lut[3935] = -9'sd11;
	qsin_lut[3936] =  9'sd0;
	icos_lut[3936] = -9'sd9;
	qsin_lut[3937] = -9'sd2;
	icos_lut[3937] = -9'sd9;
	qsin_lut[3938] = -9'sd3;
	icos_lut[3938] = -9'sd8;
	qsin_lut[3939] = -9'sd5;
	icos_lut[3939] = -9'sd7;
	qsin_lut[3940] = -9'sd6;
	icos_lut[3940] = -9'sd6;
	qsin_lut[3941] = -9'sd7;
	icos_lut[3941] = -9'sd5;
	qsin_lut[3942] = -9'sd8;
	icos_lut[3942] = -9'sd3;
	qsin_lut[3943] = -9'sd9;
	icos_lut[3943] = -9'sd2;
	qsin_lut[3944] = -9'sd9;
	icos_lut[3944] = -9'sd0;
	qsin_lut[3945] = -9'sd9;
	icos_lut[3945] =  9'sd2;
	qsin_lut[3946] = -9'sd8;
	icos_lut[3946] =  9'sd3;
	qsin_lut[3947] = -9'sd7;
	icos_lut[3947] =  9'sd5;
	qsin_lut[3948] = -9'sd6;
	icos_lut[3948] =  9'sd6;
	qsin_lut[3949] = -9'sd5;
	icos_lut[3949] =  9'sd7;
	qsin_lut[3950] = -9'sd3;
	icos_lut[3950] =  9'sd8;
	qsin_lut[3951] = -9'sd2;
	icos_lut[3951] =  9'sd9;
	qsin_lut[3952] = -9'sd0;
	icos_lut[3952] =  9'sd9;
	qsin_lut[3953] =  9'sd2;
	icos_lut[3953] =  9'sd9;
	qsin_lut[3954] =  9'sd3;
	icos_lut[3954] =  9'sd8;
	qsin_lut[3955] =  9'sd5;
	icos_lut[3955] =  9'sd7;
	qsin_lut[3956] =  9'sd6;
	icos_lut[3956] =  9'sd6;
	qsin_lut[3957] =  9'sd7;
	icos_lut[3957] =  9'sd5;
	qsin_lut[3958] =  9'sd8;
	icos_lut[3958] =  9'sd3;
	qsin_lut[3959] =  9'sd9;
	icos_lut[3959] =  9'sd2;
	qsin_lut[3960] =  9'sd9;
	icos_lut[3960] =  9'sd0;
	qsin_lut[3961] =  9'sd9;
	icos_lut[3961] = -9'sd2;
	qsin_lut[3962] =  9'sd8;
	icos_lut[3962] = -9'sd3;
	qsin_lut[3963] =  9'sd7;
	icos_lut[3963] = -9'sd5;
	qsin_lut[3964] =  9'sd6;
	icos_lut[3964] = -9'sd6;
	qsin_lut[3965] =  9'sd5;
	icos_lut[3965] = -9'sd7;
	qsin_lut[3966] =  9'sd3;
	icos_lut[3966] = -9'sd8;
	qsin_lut[3967] =  9'sd2;
	icos_lut[3967] = -9'sd9;
	qsin_lut[3968] =  9'sd0;
	icos_lut[3968] = -9'sd7;
	qsin_lut[3969] = -9'sd1;
	icos_lut[3969] = -9'sd7;
	qsin_lut[3970] = -9'sd3;
	icos_lut[3970] = -9'sd6;
	qsin_lut[3971] = -9'sd4;
	icos_lut[3971] = -9'sd6;
	qsin_lut[3972] = -9'sd5;
	icos_lut[3972] = -9'sd5;
	qsin_lut[3973] = -9'sd6;
	icos_lut[3973] = -9'sd4;
	qsin_lut[3974] = -9'sd6;
	icos_lut[3974] = -9'sd3;
	qsin_lut[3975] = -9'sd7;
	icos_lut[3975] = -9'sd1;
	qsin_lut[3976] = -9'sd7;
	icos_lut[3976] = -9'sd0;
	qsin_lut[3977] = -9'sd7;
	icos_lut[3977] =  9'sd1;
	qsin_lut[3978] = -9'sd6;
	icos_lut[3978] =  9'sd3;
	qsin_lut[3979] = -9'sd6;
	icos_lut[3979] =  9'sd4;
	qsin_lut[3980] = -9'sd5;
	icos_lut[3980] =  9'sd5;
	qsin_lut[3981] = -9'sd4;
	icos_lut[3981] =  9'sd6;
	qsin_lut[3982] = -9'sd3;
	icos_lut[3982] =  9'sd6;
	qsin_lut[3983] = -9'sd1;
	icos_lut[3983] =  9'sd7;
	qsin_lut[3984] = -9'sd0;
	icos_lut[3984] =  9'sd7;
	qsin_lut[3985] =  9'sd1;
	icos_lut[3985] =  9'sd7;
	qsin_lut[3986] =  9'sd3;
	icos_lut[3986] =  9'sd6;
	qsin_lut[3987] =  9'sd4;
	icos_lut[3987] =  9'sd6;
	qsin_lut[3988] =  9'sd5;
	icos_lut[3988] =  9'sd5;
	qsin_lut[3989] =  9'sd6;
	icos_lut[3989] =  9'sd4;
	qsin_lut[3990] =  9'sd6;
	icos_lut[3990] =  9'sd3;
	qsin_lut[3991] =  9'sd7;
	icos_lut[3991] =  9'sd1;
	qsin_lut[3992] =  9'sd7;
	icos_lut[3992] =  9'sd0;
	qsin_lut[3993] =  9'sd7;
	icos_lut[3993] = -9'sd1;
	qsin_lut[3994] =  9'sd6;
	icos_lut[3994] = -9'sd3;
	qsin_lut[3995] =  9'sd6;
	icos_lut[3995] = -9'sd4;
	qsin_lut[3996] =  9'sd5;
	icos_lut[3996] = -9'sd5;
	qsin_lut[3997] =  9'sd4;
	icos_lut[3997] = -9'sd6;
	qsin_lut[3998] =  9'sd3;
	icos_lut[3998] = -9'sd6;
	qsin_lut[3999] =  9'sd1;
	icos_lut[3999] = -9'sd7;
	qsin_lut[4000] =  9'sd0;
	icos_lut[4000] = -9'sd5;
	qsin_lut[4001] = -9'sd1;
	icos_lut[4001] = -9'sd5;
	qsin_lut[4002] = -9'sd2;
	icos_lut[4002] = -9'sd5;
	qsin_lut[4003] = -9'sd3;
	icos_lut[4003] = -9'sd4;
	qsin_lut[4004] = -9'sd4;
	icos_lut[4004] = -9'sd4;
	qsin_lut[4005] = -9'sd4;
	icos_lut[4005] = -9'sd3;
	qsin_lut[4006] = -9'sd5;
	icos_lut[4006] = -9'sd2;
	qsin_lut[4007] = -9'sd5;
	icos_lut[4007] = -9'sd1;
	qsin_lut[4008] = -9'sd5;
	icos_lut[4008] = -9'sd0;
	qsin_lut[4009] = -9'sd5;
	icos_lut[4009] =  9'sd1;
	qsin_lut[4010] = -9'sd5;
	icos_lut[4010] =  9'sd2;
	qsin_lut[4011] = -9'sd4;
	icos_lut[4011] =  9'sd3;
	qsin_lut[4012] = -9'sd4;
	icos_lut[4012] =  9'sd4;
	qsin_lut[4013] = -9'sd3;
	icos_lut[4013] =  9'sd4;
	qsin_lut[4014] = -9'sd2;
	icos_lut[4014] =  9'sd5;
	qsin_lut[4015] = -9'sd1;
	icos_lut[4015] =  9'sd5;
	qsin_lut[4016] = -9'sd0;
	icos_lut[4016] =  9'sd5;
	qsin_lut[4017] =  9'sd1;
	icos_lut[4017] =  9'sd5;
	qsin_lut[4018] =  9'sd2;
	icos_lut[4018] =  9'sd5;
	qsin_lut[4019] =  9'sd3;
	icos_lut[4019] =  9'sd4;
	qsin_lut[4020] =  9'sd4;
	icos_lut[4020] =  9'sd4;
	qsin_lut[4021] =  9'sd4;
	icos_lut[4021] =  9'sd3;
	qsin_lut[4022] =  9'sd5;
	icos_lut[4022] =  9'sd2;
	qsin_lut[4023] =  9'sd5;
	icos_lut[4023] =  9'sd1;
	qsin_lut[4024] =  9'sd5;
	icos_lut[4024] =  9'sd0;
	qsin_lut[4025] =  9'sd5;
	icos_lut[4025] = -9'sd1;
	qsin_lut[4026] =  9'sd5;
	icos_lut[4026] = -9'sd2;
	qsin_lut[4027] =  9'sd4;
	icos_lut[4027] = -9'sd3;
	qsin_lut[4028] =  9'sd4;
	icos_lut[4028] = -9'sd4;
	qsin_lut[4029] =  9'sd3;
	icos_lut[4029] = -9'sd4;
	qsin_lut[4030] =  9'sd2;
	icos_lut[4030] = -9'sd5;
	qsin_lut[4031] =  9'sd1;
	icos_lut[4031] = -9'sd5;
	qsin_lut[4032] =  9'sd0;
	icos_lut[4032] = -9'sd3;
	qsin_lut[4033] = -9'sd1;
	icos_lut[4033] = -9'sd3;
	qsin_lut[4034] = -9'sd1;
	icos_lut[4034] = -9'sd3;
	qsin_lut[4035] = -9'sd2;
	icos_lut[4035] = -9'sd2;
	qsin_lut[4036] = -9'sd2;
	icos_lut[4036] = -9'sd2;
	qsin_lut[4037] = -9'sd2;
	icos_lut[4037] = -9'sd2;
	qsin_lut[4038] = -9'sd3;
	icos_lut[4038] = -9'sd1;
	qsin_lut[4039] = -9'sd3;
	icos_lut[4039] = -9'sd1;
	qsin_lut[4040] = -9'sd3;
	icos_lut[4040] = -9'sd0;
	qsin_lut[4041] = -9'sd3;
	icos_lut[4041] =  9'sd1;
	qsin_lut[4042] = -9'sd3;
	icos_lut[4042] =  9'sd1;
	qsin_lut[4043] = -9'sd2;
	icos_lut[4043] =  9'sd2;
	qsin_lut[4044] = -9'sd2;
	icos_lut[4044] =  9'sd2;
	qsin_lut[4045] = -9'sd2;
	icos_lut[4045] =  9'sd2;
	qsin_lut[4046] = -9'sd1;
	icos_lut[4046] =  9'sd3;
	qsin_lut[4047] = -9'sd1;
	icos_lut[4047] =  9'sd3;
	qsin_lut[4048] = -9'sd0;
	icos_lut[4048] =  9'sd3;
	qsin_lut[4049] =  9'sd1;
	icos_lut[4049] =  9'sd3;
	qsin_lut[4050] =  9'sd1;
	icos_lut[4050] =  9'sd3;
	qsin_lut[4051] =  9'sd2;
	icos_lut[4051] =  9'sd2;
	qsin_lut[4052] =  9'sd2;
	icos_lut[4052] =  9'sd2;
	qsin_lut[4053] =  9'sd2;
	icos_lut[4053] =  9'sd2;
	qsin_lut[4054] =  9'sd3;
	icos_lut[4054] =  9'sd1;
	qsin_lut[4055] =  9'sd3;
	icos_lut[4055] =  9'sd1;
	qsin_lut[4056] =  9'sd3;
	icos_lut[4056] =  9'sd0;
	qsin_lut[4057] =  9'sd3;
	icos_lut[4057] = -9'sd1;
	qsin_lut[4058] =  9'sd3;
	icos_lut[4058] = -9'sd1;
	qsin_lut[4059] =  9'sd2;
	icos_lut[4059] = -9'sd2;
	qsin_lut[4060] =  9'sd2;
	icos_lut[4060] = -9'sd2;
	qsin_lut[4061] =  9'sd2;
	icos_lut[4061] = -9'sd2;
	qsin_lut[4062] =  9'sd1;
	icos_lut[4062] = -9'sd3;
	qsin_lut[4063] =  9'sd1;
	icos_lut[4063] = -9'sd3;
	qsin_lut[4064] =  9'sd0;
	icos_lut[4064] = -9'sd1;
	qsin_lut[4065] = -9'sd0;
	icos_lut[4065] = -9'sd1;
	qsin_lut[4066] = -9'sd0;
	icos_lut[4066] = -9'sd1;
	qsin_lut[4067] = -9'sd1;
	icos_lut[4067] = -9'sd1;
	qsin_lut[4068] = -9'sd1;
	icos_lut[4068] = -9'sd1;
	qsin_lut[4069] = -9'sd1;
	icos_lut[4069] = -9'sd1;
	qsin_lut[4070] = -9'sd1;
	icos_lut[4070] = -9'sd0;
	qsin_lut[4071] = -9'sd1;
	icos_lut[4071] = -9'sd0;
	qsin_lut[4072] = -9'sd1;
	icos_lut[4072] = -9'sd0;
	qsin_lut[4073] = -9'sd1;
	icos_lut[4073] =  9'sd0;
	qsin_lut[4074] = -9'sd1;
	icos_lut[4074] =  9'sd0;
	qsin_lut[4075] = -9'sd1;
	icos_lut[4075] =  9'sd1;
	qsin_lut[4076] = -9'sd1;
	icos_lut[4076] =  9'sd1;
	qsin_lut[4077] = -9'sd1;
	icos_lut[4077] =  9'sd1;
	qsin_lut[4078] = -9'sd0;
	icos_lut[4078] =  9'sd1;
	qsin_lut[4079] = -9'sd0;
	icos_lut[4079] =  9'sd1;
	qsin_lut[4080] = -9'sd0;
	icos_lut[4080] =  9'sd1;
	qsin_lut[4081] =  9'sd0;
	icos_lut[4081] =  9'sd1;
	qsin_lut[4082] =  9'sd0;
	icos_lut[4082] =  9'sd1;
	qsin_lut[4083] =  9'sd1;
	icos_lut[4083] =  9'sd1;
	qsin_lut[4084] =  9'sd1;
	icos_lut[4084] =  9'sd1;
	qsin_lut[4085] =  9'sd1;
	icos_lut[4085] =  9'sd1;
	qsin_lut[4086] =  9'sd1;
	icos_lut[4086] =  9'sd0;
	qsin_lut[4087] =  9'sd1;
	icos_lut[4087] =  9'sd0;
	qsin_lut[4088] =  9'sd1;
	icos_lut[4088] =  9'sd0;
	qsin_lut[4089] =  9'sd1;
	icos_lut[4089] = -9'sd0;
	qsin_lut[4090] =  9'sd1;
	icos_lut[4090] = -9'sd0;
	qsin_lut[4091] =  9'sd1;
	icos_lut[4091] = -9'sd1;
	qsin_lut[4092] =  9'sd1;
	icos_lut[4092] = -9'sd1;
	qsin_lut[4093] =  9'sd1;
	icos_lut[4093] = -9'sd1;
	qsin_lut[4094] =  9'sd0;
	icos_lut[4094] = -9'sd1;
	qsin_lut[4095] =  9'sd0;
	icos_lut[4095] = -9'sd1;
	qsin_lut[4096] =  9'sd0;
	icos_lut[4096] =  9'sd1;
	qsin_lut[4097] =  9'sd0;
	icos_lut[4097] =  9'sd1;
	qsin_lut[4098] =  9'sd0;
	icos_lut[4098] =  9'sd1;
	qsin_lut[4099] =  9'sd1;
	icos_lut[4099] =  9'sd1;
	qsin_lut[4100] =  9'sd1;
	icos_lut[4100] =  9'sd1;
	qsin_lut[4101] =  9'sd1;
	icos_lut[4101] =  9'sd1;
	qsin_lut[4102] =  9'sd1;
	icos_lut[4102] =  9'sd0;
	qsin_lut[4103] =  9'sd1;
	icos_lut[4103] =  9'sd0;
	qsin_lut[4104] =  9'sd1;
	icos_lut[4104] =  9'sd0;
	qsin_lut[4105] =  9'sd1;
	icos_lut[4105] = -9'sd0;
	qsin_lut[4106] =  9'sd1;
	icos_lut[4106] = -9'sd0;
	qsin_lut[4107] =  9'sd1;
	icos_lut[4107] = -9'sd1;
	qsin_lut[4108] =  9'sd1;
	icos_lut[4108] = -9'sd1;
	qsin_lut[4109] =  9'sd1;
	icos_lut[4109] = -9'sd1;
	qsin_lut[4110] =  9'sd0;
	icos_lut[4110] = -9'sd1;
	qsin_lut[4111] =  9'sd0;
	icos_lut[4111] = -9'sd1;
	qsin_lut[4112] =  9'sd0;
	icos_lut[4112] = -9'sd1;
	qsin_lut[4113] = -9'sd0;
	icos_lut[4113] = -9'sd1;
	qsin_lut[4114] = -9'sd0;
	icos_lut[4114] = -9'sd1;
	qsin_lut[4115] = -9'sd1;
	icos_lut[4115] = -9'sd1;
	qsin_lut[4116] = -9'sd1;
	icos_lut[4116] = -9'sd1;
	qsin_lut[4117] = -9'sd1;
	icos_lut[4117] = -9'sd1;
	qsin_lut[4118] = -9'sd1;
	icos_lut[4118] = -9'sd0;
	qsin_lut[4119] = -9'sd1;
	icos_lut[4119] = -9'sd0;
	qsin_lut[4120] = -9'sd1;
	icos_lut[4120] = -9'sd0;
	qsin_lut[4121] = -9'sd1;
	icos_lut[4121] =  9'sd0;
	qsin_lut[4122] = -9'sd1;
	icos_lut[4122] =  9'sd0;
	qsin_lut[4123] = -9'sd1;
	icos_lut[4123] =  9'sd1;
	qsin_lut[4124] = -9'sd1;
	icos_lut[4124] =  9'sd1;
	qsin_lut[4125] = -9'sd1;
	icos_lut[4125] =  9'sd1;
	qsin_lut[4126] = -9'sd0;
	icos_lut[4126] =  9'sd1;
	qsin_lut[4127] = -9'sd0;
	icos_lut[4127] =  9'sd1;
	qsin_lut[4128] =  9'sd0;
	icos_lut[4128] =  9'sd3;
	qsin_lut[4129] =  9'sd1;
	icos_lut[4129] =  9'sd3;
	qsin_lut[4130] =  9'sd1;
	icos_lut[4130] =  9'sd3;
	qsin_lut[4131] =  9'sd2;
	icos_lut[4131] =  9'sd2;
	qsin_lut[4132] =  9'sd2;
	icos_lut[4132] =  9'sd2;
	qsin_lut[4133] =  9'sd2;
	icos_lut[4133] =  9'sd2;
	qsin_lut[4134] =  9'sd3;
	icos_lut[4134] =  9'sd1;
	qsin_lut[4135] =  9'sd3;
	icos_lut[4135] =  9'sd1;
	qsin_lut[4136] =  9'sd3;
	icos_lut[4136] =  9'sd0;
	qsin_lut[4137] =  9'sd3;
	icos_lut[4137] = -9'sd1;
	qsin_lut[4138] =  9'sd3;
	icos_lut[4138] = -9'sd1;
	qsin_lut[4139] =  9'sd2;
	icos_lut[4139] = -9'sd2;
	qsin_lut[4140] =  9'sd2;
	icos_lut[4140] = -9'sd2;
	qsin_lut[4141] =  9'sd2;
	icos_lut[4141] = -9'sd2;
	qsin_lut[4142] =  9'sd1;
	icos_lut[4142] = -9'sd3;
	qsin_lut[4143] =  9'sd1;
	icos_lut[4143] = -9'sd3;
	qsin_lut[4144] =  9'sd0;
	icos_lut[4144] = -9'sd3;
	qsin_lut[4145] = -9'sd1;
	icos_lut[4145] = -9'sd3;
	qsin_lut[4146] = -9'sd1;
	icos_lut[4146] = -9'sd3;
	qsin_lut[4147] = -9'sd2;
	icos_lut[4147] = -9'sd2;
	qsin_lut[4148] = -9'sd2;
	icos_lut[4148] = -9'sd2;
	qsin_lut[4149] = -9'sd2;
	icos_lut[4149] = -9'sd2;
	qsin_lut[4150] = -9'sd3;
	icos_lut[4150] = -9'sd1;
	qsin_lut[4151] = -9'sd3;
	icos_lut[4151] = -9'sd1;
	qsin_lut[4152] = -9'sd3;
	icos_lut[4152] = -9'sd0;
	qsin_lut[4153] = -9'sd3;
	icos_lut[4153] =  9'sd1;
	qsin_lut[4154] = -9'sd3;
	icos_lut[4154] =  9'sd1;
	qsin_lut[4155] = -9'sd2;
	icos_lut[4155] =  9'sd2;
	qsin_lut[4156] = -9'sd2;
	icos_lut[4156] =  9'sd2;
	qsin_lut[4157] = -9'sd2;
	icos_lut[4157] =  9'sd2;
	qsin_lut[4158] = -9'sd1;
	icos_lut[4158] =  9'sd3;
	qsin_lut[4159] = -9'sd1;
	icos_lut[4159] =  9'sd3;
	qsin_lut[4160] =  9'sd0;
	icos_lut[4160] =  9'sd5;
	qsin_lut[4161] =  9'sd1;
	icos_lut[4161] =  9'sd5;
	qsin_lut[4162] =  9'sd2;
	icos_lut[4162] =  9'sd5;
	qsin_lut[4163] =  9'sd3;
	icos_lut[4163] =  9'sd4;
	qsin_lut[4164] =  9'sd4;
	icos_lut[4164] =  9'sd4;
	qsin_lut[4165] =  9'sd4;
	icos_lut[4165] =  9'sd3;
	qsin_lut[4166] =  9'sd5;
	icos_lut[4166] =  9'sd2;
	qsin_lut[4167] =  9'sd5;
	icos_lut[4167] =  9'sd1;
	qsin_lut[4168] =  9'sd5;
	icos_lut[4168] =  9'sd0;
	qsin_lut[4169] =  9'sd5;
	icos_lut[4169] = -9'sd1;
	qsin_lut[4170] =  9'sd5;
	icos_lut[4170] = -9'sd2;
	qsin_lut[4171] =  9'sd4;
	icos_lut[4171] = -9'sd3;
	qsin_lut[4172] =  9'sd4;
	icos_lut[4172] = -9'sd4;
	qsin_lut[4173] =  9'sd3;
	icos_lut[4173] = -9'sd4;
	qsin_lut[4174] =  9'sd2;
	icos_lut[4174] = -9'sd5;
	qsin_lut[4175] =  9'sd1;
	icos_lut[4175] = -9'sd5;
	qsin_lut[4176] =  9'sd0;
	icos_lut[4176] = -9'sd5;
	qsin_lut[4177] = -9'sd1;
	icos_lut[4177] = -9'sd5;
	qsin_lut[4178] = -9'sd2;
	icos_lut[4178] = -9'sd5;
	qsin_lut[4179] = -9'sd3;
	icos_lut[4179] = -9'sd4;
	qsin_lut[4180] = -9'sd4;
	icos_lut[4180] = -9'sd4;
	qsin_lut[4181] = -9'sd4;
	icos_lut[4181] = -9'sd3;
	qsin_lut[4182] = -9'sd5;
	icos_lut[4182] = -9'sd2;
	qsin_lut[4183] = -9'sd5;
	icos_lut[4183] = -9'sd1;
	qsin_lut[4184] = -9'sd5;
	icos_lut[4184] = -9'sd0;
	qsin_lut[4185] = -9'sd5;
	icos_lut[4185] =  9'sd1;
	qsin_lut[4186] = -9'sd5;
	icos_lut[4186] =  9'sd2;
	qsin_lut[4187] = -9'sd4;
	icos_lut[4187] =  9'sd3;
	qsin_lut[4188] = -9'sd4;
	icos_lut[4188] =  9'sd4;
	qsin_lut[4189] = -9'sd3;
	icos_lut[4189] =  9'sd4;
	qsin_lut[4190] = -9'sd2;
	icos_lut[4190] =  9'sd5;
	qsin_lut[4191] = -9'sd1;
	icos_lut[4191] =  9'sd5;
	qsin_lut[4192] =  9'sd0;
	icos_lut[4192] =  9'sd7;
	qsin_lut[4193] =  9'sd1;
	icos_lut[4193] =  9'sd7;
	qsin_lut[4194] =  9'sd3;
	icos_lut[4194] =  9'sd6;
	qsin_lut[4195] =  9'sd4;
	icos_lut[4195] =  9'sd6;
	qsin_lut[4196] =  9'sd5;
	icos_lut[4196] =  9'sd5;
	qsin_lut[4197] =  9'sd6;
	icos_lut[4197] =  9'sd4;
	qsin_lut[4198] =  9'sd6;
	icos_lut[4198] =  9'sd3;
	qsin_lut[4199] =  9'sd7;
	icos_lut[4199] =  9'sd1;
	qsin_lut[4200] =  9'sd7;
	icos_lut[4200] =  9'sd0;
	qsin_lut[4201] =  9'sd7;
	icos_lut[4201] = -9'sd1;
	qsin_lut[4202] =  9'sd6;
	icos_lut[4202] = -9'sd3;
	qsin_lut[4203] =  9'sd6;
	icos_lut[4203] = -9'sd4;
	qsin_lut[4204] =  9'sd5;
	icos_lut[4204] = -9'sd5;
	qsin_lut[4205] =  9'sd4;
	icos_lut[4205] = -9'sd6;
	qsin_lut[4206] =  9'sd3;
	icos_lut[4206] = -9'sd6;
	qsin_lut[4207] =  9'sd1;
	icos_lut[4207] = -9'sd7;
	qsin_lut[4208] =  9'sd0;
	icos_lut[4208] = -9'sd7;
	qsin_lut[4209] = -9'sd1;
	icos_lut[4209] = -9'sd7;
	qsin_lut[4210] = -9'sd3;
	icos_lut[4210] = -9'sd6;
	qsin_lut[4211] = -9'sd4;
	icos_lut[4211] = -9'sd6;
	qsin_lut[4212] = -9'sd5;
	icos_lut[4212] = -9'sd5;
	qsin_lut[4213] = -9'sd6;
	icos_lut[4213] = -9'sd4;
	qsin_lut[4214] = -9'sd6;
	icos_lut[4214] = -9'sd3;
	qsin_lut[4215] = -9'sd7;
	icos_lut[4215] = -9'sd1;
	qsin_lut[4216] = -9'sd7;
	icos_lut[4216] = -9'sd0;
	qsin_lut[4217] = -9'sd7;
	icos_lut[4217] =  9'sd1;
	qsin_lut[4218] = -9'sd6;
	icos_lut[4218] =  9'sd3;
	qsin_lut[4219] = -9'sd6;
	icos_lut[4219] =  9'sd4;
	qsin_lut[4220] = -9'sd5;
	icos_lut[4220] =  9'sd5;
	qsin_lut[4221] = -9'sd4;
	icos_lut[4221] =  9'sd6;
	qsin_lut[4222] = -9'sd3;
	icos_lut[4222] =  9'sd6;
	qsin_lut[4223] = -9'sd1;
	icos_lut[4223] =  9'sd7;
	qsin_lut[4224] =  9'sd0;
	icos_lut[4224] =  9'sd9;
	qsin_lut[4225] =  9'sd2;
	icos_lut[4225] =  9'sd9;
	qsin_lut[4226] =  9'sd3;
	icos_lut[4226] =  9'sd8;
	qsin_lut[4227] =  9'sd5;
	icos_lut[4227] =  9'sd7;
	qsin_lut[4228] =  9'sd6;
	icos_lut[4228] =  9'sd6;
	qsin_lut[4229] =  9'sd7;
	icos_lut[4229] =  9'sd5;
	qsin_lut[4230] =  9'sd8;
	icos_lut[4230] =  9'sd3;
	qsin_lut[4231] =  9'sd9;
	icos_lut[4231] =  9'sd2;
	qsin_lut[4232] =  9'sd9;
	icos_lut[4232] =  9'sd0;
	qsin_lut[4233] =  9'sd9;
	icos_lut[4233] = -9'sd2;
	qsin_lut[4234] =  9'sd8;
	icos_lut[4234] = -9'sd3;
	qsin_lut[4235] =  9'sd7;
	icos_lut[4235] = -9'sd5;
	qsin_lut[4236] =  9'sd6;
	icos_lut[4236] = -9'sd6;
	qsin_lut[4237] =  9'sd5;
	icos_lut[4237] = -9'sd7;
	qsin_lut[4238] =  9'sd3;
	icos_lut[4238] = -9'sd8;
	qsin_lut[4239] =  9'sd2;
	icos_lut[4239] = -9'sd9;
	qsin_lut[4240] =  9'sd0;
	icos_lut[4240] = -9'sd9;
	qsin_lut[4241] = -9'sd2;
	icos_lut[4241] = -9'sd9;
	qsin_lut[4242] = -9'sd3;
	icos_lut[4242] = -9'sd8;
	qsin_lut[4243] = -9'sd5;
	icos_lut[4243] = -9'sd7;
	qsin_lut[4244] = -9'sd6;
	icos_lut[4244] = -9'sd6;
	qsin_lut[4245] = -9'sd7;
	icos_lut[4245] = -9'sd5;
	qsin_lut[4246] = -9'sd8;
	icos_lut[4246] = -9'sd3;
	qsin_lut[4247] = -9'sd9;
	icos_lut[4247] = -9'sd2;
	qsin_lut[4248] = -9'sd9;
	icos_lut[4248] = -9'sd0;
	qsin_lut[4249] = -9'sd9;
	icos_lut[4249] =  9'sd2;
	qsin_lut[4250] = -9'sd8;
	icos_lut[4250] =  9'sd3;
	qsin_lut[4251] = -9'sd7;
	icos_lut[4251] =  9'sd5;
	qsin_lut[4252] = -9'sd6;
	icos_lut[4252] =  9'sd6;
	qsin_lut[4253] = -9'sd5;
	icos_lut[4253] =  9'sd7;
	qsin_lut[4254] = -9'sd3;
	icos_lut[4254] =  9'sd8;
	qsin_lut[4255] = -9'sd2;
	icos_lut[4255] =  9'sd9;
	qsin_lut[4256] =  9'sd0;
	icos_lut[4256] =  9'sd11;
	qsin_lut[4257] =  9'sd2;
	icos_lut[4257] =  9'sd11;
	qsin_lut[4258] =  9'sd4;
	icos_lut[4258] =  9'sd10;
	qsin_lut[4259] =  9'sd6;
	icos_lut[4259] =  9'sd9;
	qsin_lut[4260] =  9'sd8;
	icos_lut[4260] =  9'sd8;
	qsin_lut[4261] =  9'sd9;
	icos_lut[4261] =  9'sd6;
	qsin_lut[4262] =  9'sd10;
	icos_lut[4262] =  9'sd4;
	qsin_lut[4263] =  9'sd11;
	icos_lut[4263] =  9'sd2;
	qsin_lut[4264] =  9'sd11;
	icos_lut[4264] =  9'sd0;
	qsin_lut[4265] =  9'sd11;
	icos_lut[4265] = -9'sd2;
	qsin_lut[4266] =  9'sd10;
	icos_lut[4266] = -9'sd4;
	qsin_lut[4267] =  9'sd9;
	icos_lut[4267] = -9'sd6;
	qsin_lut[4268] =  9'sd8;
	icos_lut[4268] = -9'sd8;
	qsin_lut[4269] =  9'sd6;
	icos_lut[4269] = -9'sd9;
	qsin_lut[4270] =  9'sd4;
	icos_lut[4270] = -9'sd10;
	qsin_lut[4271] =  9'sd2;
	icos_lut[4271] = -9'sd11;
	qsin_lut[4272] =  9'sd0;
	icos_lut[4272] = -9'sd11;
	qsin_lut[4273] = -9'sd2;
	icos_lut[4273] = -9'sd11;
	qsin_lut[4274] = -9'sd4;
	icos_lut[4274] = -9'sd10;
	qsin_lut[4275] = -9'sd6;
	icos_lut[4275] = -9'sd9;
	qsin_lut[4276] = -9'sd8;
	icos_lut[4276] = -9'sd8;
	qsin_lut[4277] = -9'sd9;
	icos_lut[4277] = -9'sd6;
	qsin_lut[4278] = -9'sd10;
	icos_lut[4278] = -9'sd4;
	qsin_lut[4279] = -9'sd11;
	icos_lut[4279] = -9'sd2;
	qsin_lut[4280] = -9'sd11;
	icos_lut[4280] = -9'sd0;
	qsin_lut[4281] = -9'sd11;
	icos_lut[4281] =  9'sd2;
	qsin_lut[4282] = -9'sd10;
	icos_lut[4282] =  9'sd4;
	qsin_lut[4283] = -9'sd9;
	icos_lut[4283] =  9'sd6;
	qsin_lut[4284] = -9'sd8;
	icos_lut[4284] =  9'sd8;
	qsin_lut[4285] = -9'sd6;
	icos_lut[4285] =  9'sd9;
	qsin_lut[4286] = -9'sd4;
	icos_lut[4286] =  9'sd10;
	qsin_lut[4287] = -9'sd2;
	icos_lut[4287] =  9'sd11;
	qsin_lut[4288] =  9'sd0;
	icos_lut[4288] =  9'sd13;
	qsin_lut[4289] =  9'sd3;
	icos_lut[4289] =  9'sd13;
	qsin_lut[4290] =  9'sd5;
	icos_lut[4290] =  9'sd12;
	qsin_lut[4291] =  9'sd7;
	icos_lut[4291] =  9'sd11;
	qsin_lut[4292] =  9'sd9;
	icos_lut[4292] =  9'sd9;
	qsin_lut[4293] =  9'sd11;
	icos_lut[4293] =  9'sd7;
	qsin_lut[4294] =  9'sd12;
	icos_lut[4294] =  9'sd5;
	qsin_lut[4295] =  9'sd13;
	icos_lut[4295] =  9'sd3;
	qsin_lut[4296] =  9'sd13;
	icos_lut[4296] =  9'sd0;
	qsin_lut[4297] =  9'sd13;
	icos_lut[4297] = -9'sd3;
	qsin_lut[4298] =  9'sd12;
	icos_lut[4298] = -9'sd5;
	qsin_lut[4299] =  9'sd11;
	icos_lut[4299] = -9'sd7;
	qsin_lut[4300] =  9'sd9;
	icos_lut[4300] = -9'sd9;
	qsin_lut[4301] =  9'sd7;
	icos_lut[4301] = -9'sd11;
	qsin_lut[4302] =  9'sd5;
	icos_lut[4302] = -9'sd12;
	qsin_lut[4303] =  9'sd3;
	icos_lut[4303] = -9'sd13;
	qsin_lut[4304] =  9'sd0;
	icos_lut[4304] = -9'sd13;
	qsin_lut[4305] = -9'sd3;
	icos_lut[4305] = -9'sd13;
	qsin_lut[4306] = -9'sd5;
	icos_lut[4306] = -9'sd12;
	qsin_lut[4307] = -9'sd7;
	icos_lut[4307] = -9'sd11;
	qsin_lut[4308] = -9'sd9;
	icos_lut[4308] = -9'sd9;
	qsin_lut[4309] = -9'sd11;
	icos_lut[4309] = -9'sd7;
	qsin_lut[4310] = -9'sd12;
	icos_lut[4310] = -9'sd5;
	qsin_lut[4311] = -9'sd13;
	icos_lut[4311] = -9'sd3;
	qsin_lut[4312] = -9'sd13;
	icos_lut[4312] = -9'sd0;
	qsin_lut[4313] = -9'sd13;
	icos_lut[4313] =  9'sd3;
	qsin_lut[4314] = -9'sd12;
	icos_lut[4314] =  9'sd5;
	qsin_lut[4315] = -9'sd11;
	icos_lut[4315] =  9'sd7;
	qsin_lut[4316] = -9'sd9;
	icos_lut[4316] =  9'sd9;
	qsin_lut[4317] = -9'sd7;
	icos_lut[4317] =  9'sd11;
	qsin_lut[4318] = -9'sd5;
	icos_lut[4318] =  9'sd12;
	qsin_lut[4319] = -9'sd3;
	icos_lut[4319] =  9'sd13;
	qsin_lut[4320] =  9'sd0;
	icos_lut[4320] =  9'sd15;
	qsin_lut[4321] =  9'sd3;
	icos_lut[4321] =  9'sd15;
	qsin_lut[4322] =  9'sd6;
	icos_lut[4322] =  9'sd14;
	qsin_lut[4323] =  9'sd8;
	icos_lut[4323] =  9'sd12;
	qsin_lut[4324] =  9'sd11;
	icos_lut[4324] =  9'sd11;
	qsin_lut[4325] =  9'sd12;
	icos_lut[4325] =  9'sd8;
	qsin_lut[4326] =  9'sd14;
	icos_lut[4326] =  9'sd6;
	qsin_lut[4327] =  9'sd15;
	icos_lut[4327] =  9'sd3;
	qsin_lut[4328] =  9'sd15;
	icos_lut[4328] =  9'sd0;
	qsin_lut[4329] =  9'sd15;
	icos_lut[4329] = -9'sd3;
	qsin_lut[4330] =  9'sd14;
	icos_lut[4330] = -9'sd6;
	qsin_lut[4331] =  9'sd12;
	icos_lut[4331] = -9'sd8;
	qsin_lut[4332] =  9'sd11;
	icos_lut[4332] = -9'sd11;
	qsin_lut[4333] =  9'sd8;
	icos_lut[4333] = -9'sd12;
	qsin_lut[4334] =  9'sd6;
	icos_lut[4334] = -9'sd14;
	qsin_lut[4335] =  9'sd3;
	icos_lut[4335] = -9'sd15;
	qsin_lut[4336] =  9'sd0;
	icos_lut[4336] = -9'sd15;
	qsin_lut[4337] = -9'sd3;
	icos_lut[4337] = -9'sd15;
	qsin_lut[4338] = -9'sd6;
	icos_lut[4338] = -9'sd14;
	qsin_lut[4339] = -9'sd8;
	icos_lut[4339] = -9'sd12;
	qsin_lut[4340] = -9'sd11;
	icos_lut[4340] = -9'sd11;
	qsin_lut[4341] = -9'sd12;
	icos_lut[4341] = -9'sd8;
	qsin_lut[4342] = -9'sd14;
	icos_lut[4342] = -9'sd6;
	qsin_lut[4343] = -9'sd15;
	icos_lut[4343] = -9'sd3;
	qsin_lut[4344] = -9'sd15;
	icos_lut[4344] = -9'sd0;
	qsin_lut[4345] = -9'sd15;
	icos_lut[4345] =  9'sd3;
	qsin_lut[4346] = -9'sd14;
	icos_lut[4346] =  9'sd6;
	qsin_lut[4347] = -9'sd12;
	icos_lut[4347] =  9'sd8;
	qsin_lut[4348] = -9'sd11;
	icos_lut[4348] =  9'sd11;
	qsin_lut[4349] = -9'sd8;
	icos_lut[4349] =  9'sd12;
	qsin_lut[4350] = -9'sd6;
	icos_lut[4350] =  9'sd14;
	qsin_lut[4351] = -9'sd3;
	icos_lut[4351] =  9'sd15;
	qsin_lut[4352] =  9'sd0;
	icos_lut[4352] =  9'sd17;
	qsin_lut[4353] =  9'sd3;
	icos_lut[4353] =  9'sd17;
	qsin_lut[4354] =  9'sd7;
	icos_lut[4354] =  9'sd16;
	qsin_lut[4355] =  9'sd9;
	icos_lut[4355] =  9'sd14;
	qsin_lut[4356] =  9'sd12;
	icos_lut[4356] =  9'sd12;
	qsin_lut[4357] =  9'sd14;
	icos_lut[4357] =  9'sd9;
	qsin_lut[4358] =  9'sd16;
	icos_lut[4358] =  9'sd7;
	qsin_lut[4359] =  9'sd17;
	icos_lut[4359] =  9'sd3;
	qsin_lut[4360] =  9'sd17;
	icos_lut[4360] =  9'sd0;
	qsin_lut[4361] =  9'sd17;
	icos_lut[4361] = -9'sd3;
	qsin_lut[4362] =  9'sd16;
	icos_lut[4362] = -9'sd7;
	qsin_lut[4363] =  9'sd14;
	icos_lut[4363] = -9'sd9;
	qsin_lut[4364] =  9'sd12;
	icos_lut[4364] = -9'sd12;
	qsin_lut[4365] =  9'sd9;
	icos_lut[4365] = -9'sd14;
	qsin_lut[4366] =  9'sd7;
	icos_lut[4366] = -9'sd16;
	qsin_lut[4367] =  9'sd3;
	icos_lut[4367] = -9'sd17;
	qsin_lut[4368] =  9'sd0;
	icos_lut[4368] = -9'sd17;
	qsin_lut[4369] = -9'sd3;
	icos_lut[4369] = -9'sd17;
	qsin_lut[4370] = -9'sd7;
	icos_lut[4370] = -9'sd16;
	qsin_lut[4371] = -9'sd9;
	icos_lut[4371] = -9'sd14;
	qsin_lut[4372] = -9'sd12;
	icos_lut[4372] = -9'sd12;
	qsin_lut[4373] = -9'sd14;
	icos_lut[4373] = -9'sd9;
	qsin_lut[4374] = -9'sd16;
	icos_lut[4374] = -9'sd7;
	qsin_lut[4375] = -9'sd17;
	icos_lut[4375] = -9'sd3;
	qsin_lut[4376] = -9'sd17;
	icos_lut[4376] = -9'sd0;
	qsin_lut[4377] = -9'sd17;
	icos_lut[4377] =  9'sd3;
	qsin_lut[4378] = -9'sd16;
	icos_lut[4378] =  9'sd7;
	qsin_lut[4379] = -9'sd14;
	icos_lut[4379] =  9'sd9;
	qsin_lut[4380] = -9'sd12;
	icos_lut[4380] =  9'sd12;
	qsin_lut[4381] = -9'sd9;
	icos_lut[4381] =  9'sd14;
	qsin_lut[4382] = -9'sd7;
	icos_lut[4382] =  9'sd16;
	qsin_lut[4383] = -9'sd3;
	icos_lut[4383] =  9'sd17;
	qsin_lut[4384] =  9'sd0;
	icos_lut[4384] =  9'sd19;
	qsin_lut[4385] =  9'sd4;
	icos_lut[4385] =  9'sd19;
	qsin_lut[4386] =  9'sd7;
	icos_lut[4386] =  9'sd18;
	qsin_lut[4387] =  9'sd11;
	icos_lut[4387] =  9'sd16;
	qsin_lut[4388] =  9'sd13;
	icos_lut[4388] =  9'sd13;
	qsin_lut[4389] =  9'sd16;
	icos_lut[4389] =  9'sd11;
	qsin_lut[4390] =  9'sd18;
	icos_lut[4390] =  9'sd7;
	qsin_lut[4391] =  9'sd19;
	icos_lut[4391] =  9'sd4;
	qsin_lut[4392] =  9'sd19;
	icos_lut[4392] =  9'sd0;
	qsin_lut[4393] =  9'sd19;
	icos_lut[4393] = -9'sd4;
	qsin_lut[4394] =  9'sd18;
	icos_lut[4394] = -9'sd7;
	qsin_lut[4395] =  9'sd16;
	icos_lut[4395] = -9'sd11;
	qsin_lut[4396] =  9'sd13;
	icos_lut[4396] = -9'sd13;
	qsin_lut[4397] =  9'sd11;
	icos_lut[4397] = -9'sd16;
	qsin_lut[4398] =  9'sd7;
	icos_lut[4398] = -9'sd18;
	qsin_lut[4399] =  9'sd4;
	icos_lut[4399] = -9'sd19;
	qsin_lut[4400] =  9'sd0;
	icos_lut[4400] = -9'sd19;
	qsin_lut[4401] = -9'sd4;
	icos_lut[4401] = -9'sd19;
	qsin_lut[4402] = -9'sd7;
	icos_lut[4402] = -9'sd18;
	qsin_lut[4403] = -9'sd11;
	icos_lut[4403] = -9'sd16;
	qsin_lut[4404] = -9'sd13;
	icos_lut[4404] = -9'sd13;
	qsin_lut[4405] = -9'sd16;
	icos_lut[4405] = -9'sd11;
	qsin_lut[4406] = -9'sd18;
	icos_lut[4406] = -9'sd7;
	qsin_lut[4407] = -9'sd19;
	icos_lut[4407] = -9'sd4;
	qsin_lut[4408] = -9'sd19;
	icos_lut[4408] = -9'sd0;
	qsin_lut[4409] = -9'sd19;
	icos_lut[4409] =  9'sd4;
	qsin_lut[4410] = -9'sd18;
	icos_lut[4410] =  9'sd7;
	qsin_lut[4411] = -9'sd16;
	icos_lut[4411] =  9'sd11;
	qsin_lut[4412] = -9'sd13;
	icos_lut[4412] =  9'sd13;
	qsin_lut[4413] = -9'sd11;
	icos_lut[4413] =  9'sd16;
	qsin_lut[4414] = -9'sd7;
	icos_lut[4414] =  9'sd18;
	qsin_lut[4415] = -9'sd4;
	icos_lut[4415] =  9'sd19;
	qsin_lut[4416] =  9'sd0;
	icos_lut[4416] =  9'sd21;
	qsin_lut[4417] =  9'sd4;
	icos_lut[4417] =  9'sd21;
	qsin_lut[4418] =  9'sd8;
	icos_lut[4418] =  9'sd19;
	qsin_lut[4419] =  9'sd12;
	icos_lut[4419] =  9'sd17;
	qsin_lut[4420] =  9'sd15;
	icos_lut[4420] =  9'sd15;
	qsin_lut[4421] =  9'sd17;
	icos_lut[4421] =  9'sd12;
	qsin_lut[4422] =  9'sd19;
	icos_lut[4422] =  9'sd8;
	qsin_lut[4423] =  9'sd21;
	icos_lut[4423] =  9'sd4;
	qsin_lut[4424] =  9'sd21;
	icos_lut[4424] =  9'sd0;
	qsin_lut[4425] =  9'sd21;
	icos_lut[4425] = -9'sd4;
	qsin_lut[4426] =  9'sd19;
	icos_lut[4426] = -9'sd8;
	qsin_lut[4427] =  9'sd17;
	icos_lut[4427] = -9'sd12;
	qsin_lut[4428] =  9'sd15;
	icos_lut[4428] = -9'sd15;
	qsin_lut[4429] =  9'sd12;
	icos_lut[4429] = -9'sd17;
	qsin_lut[4430] =  9'sd8;
	icos_lut[4430] = -9'sd19;
	qsin_lut[4431] =  9'sd4;
	icos_lut[4431] = -9'sd21;
	qsin_lut[4432] =  9'sd0;
	icos_lut[4432] = -9'sd21;
	qsin_lut[4433] = -9'sd4;
	icos_lut[4433] = -9'sd21;
	qsin_lut[4434] = -9'sd8;
	icos_lut[4434] = -9'sd19;
	qsin_lut[4435] = -9'sd12;
	icos_lut[4435] = -9'sd17;
	qsin_lut[4436] = -9'sd15;
	icos_lut[4436] = -9'sd15;
	qsin_lut[4437] = -9'sd17;
	icos_lut[4437] = -9'sd12;
	qsin_lut[4438] = -9'sd19;
	icos_lut[4438] = -9'sd8;
	qsin_lut[4439] = -9'sd21;
	icos_lut[4439] = -9'sd4;
	qsin_lut[4440] = -9'sd21;
	icos_lut[4440] = -9'sd0;
	qsin_lut[4441] = -9'sd21;
	icos_lut[4441] =  9'sd4;
	qsin_lut[4442] = -9'sd19;
	icos_lut[4442] =  9'sd8;
	qsin_lut[4443] = -9'sd17;
	icos_lut[4443] =  9'sd12;
	qsin_lut[4444] = -9'sd15;
	icos_lut[4444] =  9'sd15;
	qsin_lut[4445] = -9'sd12;
	icos_lut[4445] =  9'sd17;
	qsin_lut[4446] = -9'sd8;
	icos_lut[4446] =  9'sd19;
	qsin_lut[4447] = -9'sd4;
	icos_lut[4447] =  9'sd21;
	qsin_lut[4448] =  9'sd0;
	icos_lut[4448] =  9'sd23;
	qsin_lut[4449] =  9'sd4;
	icos_lut[4449] =  9'sd23;
	qsin_lut[4450] =  9'sd9;
	icos_lut[4450] =  9'sd21;
	qsin_lut[4451] =  9'sd13;
	icos_lut[4451] =  9'sd19;
	qsin_lut[4452] =  9'sd16;
	icos_lut[4452] =  9'sd16;
	qsin_lut[4453] =  9'sd19;
	icos_lut[4453] =  9'sd13;
	qsin_lut[4454] =  9'sd21;
	icos_lut[4454] =  9'sd9;
	qsin_lut[4455] =  9'sd23;
	icos_lut[4455] =  9'sd4;
	qsin_lut[4456] =  9'sd23;
	icos_lut[4456] =  9'sd0;
	qsin_lut[4457] =  9'sd23;
	icos_lut[4457] = -9'sd4;
	qsin_lut[4458] =  9'sd21;
	icos_lut[4458] = -9'sd9;
	qsin_lut[4459] =  9'sd19;
	icos_lut[4459] = -9'sd13;
	qsin_lut[4460] =  9'sd16;
	icos_lut[4460] = -9'sd16;
	qsin_lut[4461] =  9'sd13;
	icos_lut[4461] = -9'sd19;
	qsin_lut[4462] =  9'sd9;
	icos_lut[4462] = -9'sd21;
	qsin_lut[4463] =  9'sd4;
	icos_lut[4463] = -9'sd23;
	qsin_lut[4464] =  9'sd0;
	icos_lut[4464] = -9'sd23;
	qsin_lut[4465] = -9'sd4;
	icos_lut[4465] = -9'sd23;
	qsin_lut[4466] = -9'sd9;
	icos_lut[4466] = -9'sd21;
	qsin_lut[4467] = -9'sd13;
	icos_lut[4467] = -9'sd19;
	qsin_lut[4468] = -9'sd16;
	icos_lut[4468] = -9'sd16;
	qsin_lut[4469] = -9'sd19;
	icos_lut[4469] = -9'sd13;
	qsin_lut[4470] = -9'sd21;
	icos_lut[4470] = -9'sd9;
	qsin_lut[4471] = -9'sd23;
	icos_lut[4471] = -9'sd4;
	qsin_lut[4472] = -9'sd23;
	icos_lut[4472] = -9'sd0;
	qsin_lut[4473] = -9'sd23;
	icos_lut[4473] =  9'sd4;
	qsin_lut[4474] = -9'sd21;
	icos_lut[4474] =  9'sd9;
	qsin_lut[4475] = -9'sd19;
	icos_lut[4475] =  9'sd13;
	qsin_lut[4476] = -9'sd16;
	icos_lut[4476] =  9'sd16;
	qsin_lut[4477] = -9'sd13;
	icos_lut[4477] =  9'sd19;
	qsin_lut[4478] = -9'sd9;
	icos_lut[4478] =  9'sd21;
	qsin_lut[4479] = -9'sd4;
	icos_lut[4479] =  9'sd23;
	qsin_lut[4480] =  9'sd0;
	icos_lut[4480] =  9'sd25;
	qsin_lut[4481] =  9'sd5;
	icos_lut[4481] =  9'sd25;
	qsin_lut[4482] =  9'sd10;
	icos_lut[4482] =  9'sd23;
	qsin_lut[4483] =  9'sd14;
	icos_lut[4483] =  9'sd21;
	qsin_lut[4484] =  9'sd18;
	icos_lut[4484] =  9'sd18;
	qsin_lut[4485] =  9'sd21;
	icos_lut[4485] =  9'sd14;
	qsin_lut[4486] =  9'sd23;
	icos_lut[4486] =  9'sd10;
	qsin_lut[4487] =  9'sd25;
	icos_lut[4487] =  9'sd5;
	qsin_lut[4488] =  9'sd25;
	icos_lut[4488] =  9'sd0;
	qsin_lut[4489] =  9'sd25;
	icos_lut[4489] = -9'sd5;
	qsin_lut[4490] =  9'sd23;
	icos_lut[4490] = -9'sd10;
	qsin_lut[4491] =  9'sd21;
	icos_lut[4491] = -9'sd14;
	qsin_lut[4492] =  9'sd18;
	icos_lut[4492] = -9'sd18;
	qsin_lut[4493] =  9'sd14;
	icos_lut[4493] = -9'sd21;
	qsin_lut[4494] =  9'sd10;
	icos_lut[4494] = -9'sd23;
	qsin_lut[4495] =  9'sd5;
	icos_lut[4495] = -9'sd25;
	qsin_lut[4496] =  9'sd0;
	icos_lut[4496] = -9'sd25;
	qsin_lut[4497] = -9'sd5;
	icos_lut[4497] = -9'sd25;
	qsin_lut[4498] = -9'sd10;
	icos_lut[4498] = -9'sd23;
	qsin_lut[4499] = -9'sd14;
	icos_lut[4499] = -9'sd21;
	qsin_lut[4500] = -9'sd18;
	icos_lut[4500] = -9'sd18;
	qsin_lut[4501] = -9'sd21;
	icos_lut[4501] = -9'sd14;
	qsin_lut[4502] = -9'sd23;
	icos_lut[4502] = -9'sd10;
	qsin_lut[4503] = -9'sd25;
	icos_lut[4503] = -9'sd5;
	qsin_lut[4504] = -9'sd25;
	icos_lut[4504] = -9'sd0;
	qsin_lut[4505] = -9'sd25;
	icos_lut[4505] =  9'sd5;
	qsin_lut[4506] = -9'sd23;
	icos_lut[4506] =  9'sd10;
	qsin_lut[4507] = -9'sd21;
	icos_lut[4507] =  9'sd14;
	qsin_lut[4508] = -9'sd18;
	icos_lut[4508] =  9'sd18;
	qsin_lut[4509] = -9'sd14;
	icos_lut[4509] =  9'sd21;
	qsin_lut[4510] = -9'sd10;
	icos_lut[4510] =  9'sd23;
	qsin_lut[4511] = -9'sd5;
	icos_lut[4511] =  9'sd25;
	qsin_lut[4512] =  9'sd0;
	icos_lut[4512] =  9'sd27;
	qsin_lut[4513] =  9'sd5;
	icos_lut[4513] =  9'sd26;
	qsin_lut[4514] =  9'sd10;
	icos_lut[4514] =  9'sd25;
	qsin_lut[4515] =  9'sd15;
	icos_lut[4515] =  9'sd22;
	qsin_lut[4516] =  9'sd19;
	icos_lut[4516] =  9'sd19;
	qsin_lut[4517] =  9'sd22;
	icos_lut[4517] =  9'sd15;
	qsin_lut[4518] =  9'sd25;
	icos_lut[4518] =  9'sd10;
	qsin_lut[4519] =  9'sd26;
	icos_lut[4519] =  9'sd5;
	qsin_lut[4520] =  9'sd27;
	icos_lut[4520] =  9'sd0;
	qsin_lut[4521] =  9'sd26;
	icos_lut[4521] = -9'sd5;
	qsin_lut[4522] =  9'sd25;
	icos_lut[4522] = -9'sd10;
	qsin_lut[4523] =  9'sd22;
	icos_lut[4523] = -9'sd15;
	qsin_lut[4524] =  9'sd19;
	icos_lut[4524] = -9'sd19;
	qsin_lut[4525] =  9'sd15;
	icos_lut[4525] = -9'sd22;
	qsin_lut[4526] =  9'sd10;
	icos_lut[4526] = -9'sd25;
	qsin_lut[4527] =  9'sd5;
	icos_lut[4527] = -9'sd26;
	qsin_lut[4528] =  9'sd0;
	icos_lut[4528] = -9'sd27;
	qsin_lut[4529] = -9'sd5;
	icos_lut[4529] = -9'sd26;
	qsin_lut[4530] = -9'sd10;
	icos_lut[4530] = -9'sd25;
	qsin_lut[4531] = -9'sd15;
	icos_lut[4531] = -9'sd22;
	qsin_lut[4532] = -9'sd19;
	icos_lut[4532] = -9'sd19;
	qsin_lut[4533] = -9'sd22;
	icos_lut[4533] = -9'sd15;
	qsin_lut[4534] = -9'sd25;
	icos_lut[4534] = -9'sd10;
	qsin_lut[4535] = -9'sd26;
	icos_lut[4535] = -9'sd5;
	qsin_lut[4536] = -9'sd27;
	icos_lut[4536] = -9'sd0;
	qsin_lut[4537] = -9'sd26;
	icos_lut[4537] =  9'sd5;
	qsin_lut[4538] = -9'sd25;
	icos_lut[4538] =  9'sd10;
	qsin_lut[4539] = -9'sd22;
	icos_lut[4539] =  9'sd15;
	qsin_lut[4540] = -9'sd19;
	icos_lut[4540] =  9'sd19;
	qsin_lut[4541] = -9'sd15;
	icos_lut[4541] =  9'sd22;
	qsin_lut[4542] = -9'sd10;
	icos_lut[4542] =  9'sd25;
	qsin_lut[4543] = -9'sd5;
	icos_lut[4543] =  9'sd26;
	qsin_lut[4544] =  9'sd0;
	icos_lut[4544] =  9'sd29;
	qsin_lut[4545] =  9'sd6;
	icos_lut[4545] =  9'sd28;
	qsin_lut[4546] =  9'sd11;
	icos_lut[4546] =  9'sd27;
	qsin_lut[4547] =  9'sd16;
	icos_lut[4547] =  9'sd24;
	qsin_lut[4548] =  9'sd21;
	icos_lut[4548] =  9'sd21;
	qsin_lut[4549] =  9'sd24;
	icos_lut[4549] =  9'sd16;
	qsin_lut[4550] =  9'sd27;
	icos_lut[4550] =  9'sd11;
	qsin_lut[4551] =  9'sd28;
	icos_lut[4551] =  9'sd6;
	qsin_lut[4552] =  9'sd29;
	icos_lut[4552] =  9'sd0;
	qsin_lut[4553] =  9'sd28;
	icos_lut[4553] = -9'sd6;
	qsin_lut[4554] =  9'sd27;
	icos_lut[4554] = -9'sd11;
	qsin_lut[4555] =  9'sd24;
	icos_lut[4555] = -9'sd16;
	qsin_lut[4556] =  9'sd21;
	icos_lut[4556] = -9'sd21;
	qsin_lut[4557] =  9'sd16;
	icos_lut[4557] = -9'sd24;
	qsin_lut[4558] =  9'sd11;
	icos_lut[4558] = -9'sd27;
	qsin_lut[4559] =  9'sd6;
	icos_lut[4559] = -9'sd28;
	qsin_lut[4560] =  9'sd0;
	icos_lut[4560] = -9'sd29;
	qsin_lut[4561] = -9'sd6;
	icos_lut[4561] = -9'sd28;
	qsin_lut[4562] = -9'sd11;
	icos_lut[4562] = -9'sd27;
	qsin_lut[4563] = -9'sd16;
	icos_lut[4563] = -9'sd24;
	qsin_lut[4564] = -9'sd21;
	icos_lut[4564] = -9'sd21;
	qsin_lut[4565] = -9'sd24;
	icos_lut[4565] = -9'sd16;
	qsin_lut[4566] = -9'sd27;
	icos_lut[4566] = -9'sd11;
	qsin_lut[4567] = -9'sd28;
	icos_lut[4567] = -9'sd6;
	qsin_lut[4568] = -9'sd29;
	icos_lut[4568] = -9'sd0;
	qsin_lut[4569] = -9'sd28;
	icos_lut[4569] =  9'sd6;
	qsin_lut[4570] = -9'sd27;
	icos_lut[4570] =  9'sd11;
	qsin_lut[4571] = -9'sd24;
	icos_lut[4571] =  9'sd16;
	qsin_lut[4572] = -9'sd21;
	icos_lut[4572] =  9'sd21;
	qsin_lut[4573] = -9'sd16;
	icos_lut[4573] =  9'sd24;
	qsin_lut[4574] = -9'sd11;
	icos_lut[4574] =  9'sd27;
	qsin_lut[4575] = -9'sd6;
	icos_lut[4575] =  9'sd28;
	qsin_lut[4576] =  9'sd0;
	icos_lut[4576] =  9'sd31;
	qsin_lut[4577] =  9'sd6;
	icos_lut[4577] =  9'sd30;
	qsin_lut[4578] =  9'sd12;
	icos_lut[4578] =  9'sd29;
	qsin_lut[4579] =  9'sd17;
	icos_lut[4579] =  9'sd26;
	qsin_lut[4580] =  9'sd22;
	icos_lut[4580] =  9'sd22;
	qsin_lut[4581] =  9'sd26;
	icos_lut[4581] =  9'sd17;
	qsin_lut[4582] =  9'sd29;
	icos_lut[4582] =  9'sd12;
	qsin_lut[4583] =  9'sd30;
	icos_lut[4583] =  9'sd6;
	qsin_lut[4584] =  9'sd31;
	icos_lut[4584] =  9'sd0;
	qsin_lut[4585] =  9'sd30;
	icos_lut[4585] = -9'sd6;
	qsin_lut[4586] =  9'sd29;
	icos_lut[4586] = -9'sd12;
	qsin_lut[4587] =  9'sd26;
	icos_lut[4587] = -9'sd17;
	qsin_lut[4588] =  9'sd22;
	icos_lut[4588] = -9'sd22;
	qsin_lut[4589] =  9'sd17;
	icos_lut[4589] = -9'sd26;
	qsin_lut[4590] =  9'sd12;
	icos_lut[4590] = -9'sd29;
	qsin_lut[4591] =  9'sd6;
	icos_lut[4591] = -9'sd30;
	qsin_lut[4592] =  9'sd0;
	icos_lut[4592] = -9'sd31;
	qsin_lut[4593] = -9'sd6;
	icos_lut[4593] = -9'sd30;
	qsin_lut[4594] = -9'sd12;
	icos_lut[4594] = -9'sd29;
	qsin_lut[4595] = -9'sd17;
	icos_lut[4595] = -9'sd26;
	qsin_lut[4596] = -9'sd22;
	icos_lut[4596] = -9'sd22;
	qsin_lut[4597] = -9'sd26;
	icos_lut[4597] = -9'sd17;
	qsin_lut[4598] = -9'sd29;
	icos_lut[4598] = -9'sd12;
	qsin_lut[4599] = -9'sd30;
	icos_lut[4599] = -9'sd6;
	qsin_lut[4600] = -9'sd31;
	icos_lut[4600] = -9'sd0;
	qsin_lut[4601] = -9'sd30;
	icos_lut[4601] =  9'sd6;
	qsin_lut[4602] = -9'sd29;
	icos_lut[4602] =  9'sd12;
	qsin_lut[4603] = -9'sd26;
	icos_lut[4603] =  9'sd17;
	qsin_lut[4604] = -9'sd22;
	icos_lut[4604] =  9'sd22;
	qsin_lut[4605] = -9'sd17;
	icos_lut[4605] =  9'sd26;
	qsin_lut[4606] = -9'sd12;
	icos_lut[4606] =  9'sd29;
	qsin_lut[4607] = -9'sd6;
	icos_lut[4607] =  9'sd30;
	qsin_lut[4608] =  9'sd0;
	icos_lut[4608] =  9'sd33;
	qsin_lut[4609] =  9'sd6;
	icos_lut[4609] =  9'sd32;
	qsin_lut[4610] =  9'sd13;
	icos_lut[4610] =  9'sd30;
	qsin_lut[4611] =  9'sd18;
	icos_lut[4611] =  9'sd27;
	qsin_lut[4612] =  9'sd23;
	icos_lut[4612] =  9'sd23;
	qsin_lut[4613] =  9'sd27;
	icos_lut[4613] =  9'sd18;
	qsin_lut[4614] =  9'sd30;
	icos_lut[4614] =  9'sd13;
	qsin_lut[4615] =  9'sd32;
	icos_lut[4615] =  9'sd6;
	qsin_lut[4616] =  9'sd33;
	icos_lut[4616] =  9'sd0;
	qsin_lut[4617] =  9'sd32;
	icos_lut[4617] = -9'sd6;
	qsin_lut[4618] =  9'sd30;
	icos_lut[4618] = -9'sd13;
	qsin_lut[4619] =  9'sd27;
	icos_lut[4619] = -9'sd18;
	qsin_lut[4620] =  9'sd23;
	icos_lut[4620] = -9'sd23;
	qsin_lut[4621] =  9'sd18;
	icos_lut[4621] = -9'sd27;
	qsin_lut[4622] =  9'sd13;
	icos_lut[4622] = -9'sd30;
	qsin_lut[4623] =  9'sd6;
	icos_lut[4623] = -9'sd32;
	qsin_lut[4624] =  9'sd0;
	icos_lut[4624] = -9'sd33;
	qsin_lut[4625] = -9'sd6;
	icos_lut[4625] = -9'sd32;
	qsin_lut[4626] = -9'sd13;
	icos_lut[4626] = -9'sd30;
	qsin_lut[4627] = -9'sd18;
	icos_lut[4627] = -9'sd27;
	qsin_lut[4628] = -9'sd23;
	icos_lut[4628] = -9'sd23;
	qsin_lut[4629] = -9'sd27;
	icos_lut[4629] = -9'sd18;
	qsin_lut[4630] = -9'sd30;
	icos_lut[4630] = -9'sd13;
	qsin_lut[4631] = -9'sd32;
	icos_lut[4631] = -9'sd6;
	qsin_lut[4632] = -9'sd33;
	icos_lut[4632] = -9'sd0;
	qsin_lut[4633] = -9'sd32;
	icos_lut[4633] =  9'sd6;
	qsin_lut[4634] = -9'sd30;
	icos_lut[4634] =  9'sd13;
	qsin_lut[4635] = -9'sd27;
	icos_lut[4635] =  9'sd18;
	qsin_lut[4636] = -9'sd23;
	icos_lut[4636] =  9'sd23;
	qsin_lut[4637] = -9'sd18;
	icos_lut[4637] =  9'sd27;
	qsin_lut[4638] = -9'sd13;
	icos_lut[4638] =  9'sd30;
	qsin_lut[4639] = -9'sd6;
	icos_lut[4639] =  9'sd32;
	qsin_lut[4640] =  9'sd0;
	icos_lut[4640] =  9'sd35;
	qsin_lut[4641] =  9'sd7;
	icos_lut[4641] =  9'sd34;
	qsin_lut[4642] =  9'sd13;
	icos_lut[4642] =  9'sd32;
	qsin_lut[4643] =  9'sd19;
	icos_lut[4643] =  9'sd29;
	qsin_lut[4644] =  9'sd25;
	icos_lut[4644] =  9'sd25;
	qsin_lut[4645] =  9'sd29;
	icos_lut[4645] =  9'sd19;
	qsin_lut[4646] =  9'sd32;
	icos_lut[4646] =  9'sd13;
	qsin_lut[4647] =  9'sd34;
	icos_lut[4647] =  9'sd7;
	qsin_lut[4648] =  9'sd35;
	icos_lut[4648] =  9'sd0;
	qsin_lut[4649] =  9'sd34;
	icos_lut[4649] = -9'sd7;
	qsin_lut[4650] =  9'sd32;
	icos_lut[4650] = -9'sd13;
	qsin_lut[4651] =  9'sd29;
	icos_lut[4651] = -9'sd19;
	qsin_lut[4652] =  9'sd25;
	icos_lut[4652] = -9'sd25;
	qsin_lut[4653] =  9'sd19;
	icos_lut[4653] = -9'sd29;
	qsin_lut[4654] =  9'sd13;
	icos_lut[4654] = -9'sd32;
	qsin_lut[4655] =  9'sd7;
	icos_lut[4655] = -9'sd34;
	qsin_lut[4656] =  9'sd0;
	icos_lut[4656] = -9'sd35;
	qsin_lut[4657] = -9'sd7;
	icos_lut[4657] = -9'sd34;
	qsin_lut[4658] = -9'sd13;
	icos_lut[4658] = -9'sd32;
	qsin_lut[4659] = -9'sd19;
	icos_lut[4659] = -9'sd29;
	qsin_lut[4660] = -9'sd25;
	icos_lut[4660] = -9'sd25;
	qsin_lut[4661] = -9'sd29;
	icos_lut[4661] = -9'sd19;
	qsin_lut[4662] = -9'sd32;
	icos_lut[4662] = -9'sd13;
	qsin_lut[4663] = -9'sd34;
	icos_lut[4663] = -9'sd7;
	qsin_lut[4664] = -9'sd35;
	icos_lut[4664] = -9'sd0;
	qsin_lut[4665] = -9'sd34;
	icos_lut[4665] =  9'sd7;
	qsin_lut[4666] = -9'sd32;
	icos_lut[4666] =  9'sd13;
	qsin_lut[4667] = -9'sd29;
	icos_lut[4667] =  9'sd19;
	qsin_lut[4668] = -9'sd25;
	icos_lut[4668] =  9'sd25;
	qsin_lut[4669] = -9'sd19;
	icos_lut[4669] =  9'sd29;
	qsin_lut[4670] = -9'sd13;
	icos_lut[4670] =  9'sd32;
	qsin_lut[4671] = -9'sd7;
	icos_lut[4671] =  9'sd34;
	qsin_lut[4672] =  9'sd0;
	icos_lut[4672] =  9'sd37;
	qsin_lut[4673] =  9'sd7;
	icos_lut[4673] =  9'sd36;
	qsin_lut[4674] =  9'sd14;
	icos_lut[4674] =  9'sd34;
	qsin_lut[4675] =  9'sd21;
	icos_lut[4675] =  9'sd31;
	qsin_lut[4676] =  9'sd26;
	icos_lut[4676] =  9'sd26;
	qsin_lut[4677] =  9'sd31;
	icos_lut[4677] =  9'sd21;
	qsin_lut[4678] =  9'sd34;
	icos_lut[4678] =  9'sd14;
	qsin_lut[4679] =  9'sd36;
	icos_lut[4679] =  9'sd7;
	qsin_lut[4680] =  9'sd37;
	icos_lut[4680] =  9'sd0;
	qsin_lut[4681] =  9'sd36;
	icos_lut[4681] = -9'sd7;
	qsin_lut[4682] =  9'sd34;
	icos_lut[4682] = -9'sd14;
	qsin_lut[4683] =  9'sd31;
	icos_lut[4683] = -9'sd21;
	qsin_lut[4684] =  9'sd26;
	icos_lut[4684] = -9'sd26;
	qsin_lut[4685] =  9'sd21;
	icos_lut[4685] = -9'sd31;
	qsin_lut[4686] =  9'sd14;
	icos_lut[4686] = -9'sd34;
	qsin_lut[4687] =  9'sd7;
	icos_lut[4687] = -9'sd36;
	qsin_lut[4688] =  9'sd0;
	icos_lut[4688] = -9'sd37;
	qsin_lut[4689] = -9'sd7;
	icos_lut[4689] = -9'sd36;
	qsin_lut[4690] = -9'sd14;
	icos_lut[4690] = -9'sd34;
	qsin_lut[4691] = -9'sd21;
	icos_lut[4691] = -9'sd31;
	qsin_lut[4692] = -9'sd26;
	icos_lut[4692] = -9'sd26;
	qsin_lut[4693] = -9'sd31;
	icos_lut[4693] = -9'sd21;
	qsin_lut[4694] = -9'sd34;
	icos_lut[4694] = -9'sd14;
	qsin_lut[4695] = -9'sd36;
	icos_lut[4695] = -9'sd7;
	qsin_lut[4696] = -9'sd37;
	icos_lut[4696] = -9'sd0;
	qsin_lut[4697] = -9'sd36;
	icos_lut[4697] =  9'sd7;
	qsin_lut[4698] = -9'sd34;
	icos_lut[4698] =  9'sd14;
	qsin_lut[4699] = -9'sd31;
	icos_lut[4699] =  9'sd21;
	qsin_lut[4700] = -9'sd26;
	icos_lut[4700] =  9'sd26;
	qsin_lut[4701] = -9'sd21;
	icos_lut[4701] =  9'sd31;
	qsin_lut[4702] = -9'sd14;
	icos_lut[4702] =  9'sd34;
	qsin_lut[4703] = -9'sd7;
	icos_lut[4703] =  9'sd36;
	qsin_lut[4704] =  9'sd0;
	icos_lut[4704] =  9'sd39;
	qsin_lut[4705] =  9'sd8;
	icos_lut[4705] =  9'sd38;
	qsin_lut[4706] =  9'sd15;
	icos_lut[4706] =  9'sd36;
	qsin_lut[4707] =  9'sd22;
	icos_lut[4707] =  9'sd32;
	qsin_lut[4708] =  9'sd28;
	icos_lut[4708] =  9'sd28;
	qsin_lut[4709] =  9'sd32;
	icos_lut[4709] =  9'sd22;
	qsin_lut[4710] =  9'sd36;
	icos_lut[4710] =  9'sd15;
	qsin_lut[4711] =  9'sd38;
	icos_lut[4711] =  9'sd8;
	qsin_lut[4712] =  9'sd39;
	icos_lut[4712] =  9'sd0;
	qsin_lut[4713] =  9'sd38;
	icos_lut[4713] = -9'sd8;
	qsin_lut[4714] =  9'sd36;
	icos_lut[4714] = -9'sd15;
	qsin_lut[4715] =  9'sd32;
	icos_lut[4715] = -9'sd22;
	qsin_lut[4716] =  9'sd28;
	icos_lut[4716] = -9'sd28;
	qsin_lut[4717] =  9'sd22;
	icos_lut[4717] = -9'sd32;
	qsin_lut[4718] =  9'sd15;
	icos_lut[4718] = -9'sd36;
	qsin_lut[4719] =  9'sd8;
	icos_lut[4719] = -9'sd38;
	qsin_lut[4720] =  9'sd0;
	icos_lut[4720] = -9'sd39;
	qsin_lut[4721] = -9'sd8;
	icos_lut[4721] = -9'sd38;
	qsin_lut[4722] = -9'sd15;
	icos_lut[4722] = -9'sd36;
	qsin_lut[4723] = -9'sd22;
	icos_lut[4723] = -9'sd32;
	qsin_lut[4724] = -9'sd28;
	icos_lut[4724] = -9'sd28;
	qsin_lut[4725] = -9'sd32;
	icos_lut[4725] = -9'sd22;
	qsin_lut[4726] = -9'sd36;
	icos_lut[4726] = -9'sd15;
	qsin_lut[4727] = -9'sd38;
	icos_lut[4727] = -9'sd8;
	qsin_lut[4728] = -9'sd39;
	icos_lut[4728] = -9'sd0;
	qsin_lut[4729] = -9'sd38;
	icos_lut[4729] =  9'sd8;
	qsin_lut[4730] = -9'sd36;
	icos_lut[4730] =  9'sd15;
	qsin_lut[4731] = -9'sd32;
	icos_lut[4731] =  9'sd22;
	qsin_lut[4732] = -9'sd28;
	icos_lut[4732] =  9'sd28;
	qsin_lut[4733] = -9'sd22;
	icos_lut[4733] =  9'sd32;
	qsin_lut[4734] = -9'sd15;
	icos_lut[4734] =  9'sd36;
	qsin_lut[4735] = -9'sd8;
	icos_lut[4735] =  9'sd38;
	qsin_lut[4736] =  9'sd0;
	icos_lut[4736] =  9'sd41;
	qsin_lut[4737] =  9'sd8;
	icos_lut[4737] =  9'sd40;
	qsin_lut[4738] =  9'sd16;
	icos_lut[4738] =  9'sd38;
	qsin_lut[4739] =  9'sd23;
	icos_lut[4739] =  9'sd34;
	qsin_lut[4740] =  9'sd29;
	icos_lut[4740] =  9'sd29;
	qsin_lut[4741] =  9'sd34;
	icos_lut[4741] =  9'sd23;
	qsin_lut[4742] =  9'sd38;
	icos_lut[4742] =  9'sd16;
	qsin_lut[4743] =  9'sd40;
	icos_lut[4743] =  9'sd8;
	qsin_lut[4744] =  9'sd41;
	icos_lut[4744] =  9'sd0;
	qsin_lut[4745] =  9'sd40;
	icos_lut[4745] = -9'sd8;
	qsin_lut[4746] =  9'sd38;
	icos_lut[4746] = -9'sd16;
	qsin_lut[4747] =  9'sd34;
	icos_lut[4747] = -9'sd23;
	qsin_lut[4748] =  9'sd29;
	icos_lut[4748] = -9'sd29;
	qsin_lut[4749] =  9'sd23;
	icos_lut[4749] = -9'sd34;
	qsin_lut[4750] =  9'sd16;
	icos_lut[4750] = -9'sd38;
	qsin_lut[4751] =  9'sd8;
	icos_lut[4751] = -9'sd40;
	qsin_lut[4752] =  9'sd0;
	icos_lut[4752] = -9'sd41;
	qsin_lut[4753] = -9'sd8;
	icos_lut[4753] = -9'sd40;
	qsin_lut[4754] = -9'sd16;
	icos_lut[4754] = -9'sd38;
	qsin_lut[4755] = -9'sd23;
	icos_lut[4755] = -9'sd34;
	qsin_lut[4756] = -9'sd29;
	icos_lut[4756] = -9'sd29;
	qsin_lut[4757] = -9'sd34;
	icos_lut[4757] = -9'sd23;
	qsin_lut[4758] = -9'sd38;
	icos_lut[4758] = -9'sd16;
	qsin_lut[4759] = -9'sd40;
	icos_lut[4759] = -9'sd8;
	qsin_lut[4760] = -9'sd41;
	icos_lut[4760] = -9'sd0;
	qsin_lut[4761] = -9'sd40;
	icos_lut[4761] =  9'sd8;
	qsin_lut[4762] = -9'sd38;
	icos_lut[4762] =  9'sd16;
	qsin_lut[4763] = -9'sd34;
	icos_lut[4763] =  9'sd23;
	qsin_lut[4764] = -9'sd29;
	icos_lut[4764] =  9'sd29;
	qsin_lut[4765] = -9'sd23;
	icos_lut[4765] =  9'sd34;
	qsin_lut[4766] = -9'sd16;
	icos_lut[4766] =  9'sd38;
	qsin_lut[4767] = -9'sd8;
	icos_lut[4767] =  9'sd40;
	qsin_lut[4768] =  9'sd0;
	icos_lut[4768] =  9'sd43;
	qsin_lut[4769] =  9'sd8;
	icos_lut[4769] =  9'sd42;
	qsin_lut[4770] =  9'sd16;
	icos_lut[4770] =  9'sd40;
	qsin_lut[4771] =  9'sd24;
	icos_lut[4771] =  9'sd36;
	qsin_lut[4772] =  9'sd30;
	icos_lut[4772] =  9'sd30;
	qsin_lut[4773] =  9'sd36;
	icos_lut[4773] =  9'sd24;
	qsin_lut[4774] =  9'sd40;
	icos_lut[4774] =  9'sd16;
	qsin_lut[4775] =  9'sd42;
	icos_lut[4775] =  9'sd8;
	qsin_lut[4776] =  9'sd43;
	icos_lut[4776] =  9'sd0;
	qsin_lut[4777] =  9'sd42;
	icos_lut[4777] = -9'sd8;
	qsin_lut[4778] =  9'sd40;
	icos_lut[4778] = -9'sd16;
	qsin_lut[4779] =  9'sd36;
	icos_lut[4779] = -9'sd24;
	qsin_lut[4780] =  9'sd30;
	icos_lut[4780] = -9'sd30;
	qsin_lut[4781] =  9'sd24;
	icos_lut[4781] = -9'sd36;
	qsin_lut[4782] =  9'sd16;
	icos_lut[4782] = -9'sd40;
	qsin_lut[4783] =  9'sd8;
	icos_lut[4783] = -9'sd42;
	qsin_lut[4784] =  9'sd0;
	icos_lut[4784] = -9'sd43;
	qsin_lut[4785] = -9'sd8;
	icos_lut[4785] = -9'sd42;
	qsin_lut[4786] = -9'sd16;
	icos_lut[4786] = -9'sd40;
	qsin_lut[4787] = -9'sd24;
	icos_lut[4787] = -9'sd36;
	qsin_lut[4788] = -9'sd30;
	icos_lut[4788] = -9'sd30;
	qsin_lut[4789] = -9'sd36;
	icos_lut[4789] = -9'sd24;
	qsin_lut[4790] = -9'sd40;
	icos_lut[4790] = -9'sd16;
	qsin_lut[4791] = -9'sd42;
	icos_lut[4791] = -9'sd8;
	qsin_lut[4792] = -9'sd43;
	icos_lut[4792] = -9'sd0;
	qsin_lut[4793] = -9'sd42;
	icos_lut[4793] =  9'sd8;
	qsin_lut[4794] = -9'sd40;
	icos_lut[4794] =  9'sd16;
	qsin_lut[4795] = -9'sd36;
	icos_lut[4795] =  9'sd24;
	qsin_lut[4796] = -9'sd30;
	icos_lut[4796] =  9'sd30;
	qsin_lut[4797] = -9'sd24;
	icos_lut[4797] =  9'sd36;
	qsin_lut[4798] = -9'sd16;
	icos_lut[4798] =  9'sd40;
	qsin_lut[4799] = -9'sd8;
	icos_lut[4799] =  9'sd42;
	qsin_lut[4800] =  9'sd0;
	icos_lut[4800] =  9'sd45;
	qsin_lut[4801] =  9'sd9;
	icos_lut[4801] =  9'sd44;
	qsin_lut[4802] =  9'sd17;
	icos_lut[4802] =  9'sd42;
	qsin_lut[4803] =  9'sd25;
	icos_lut[4803] =  9'sd37;
	qsin_lut[4804] =  9'sd32;
	icos_lut[4804] =  9'sd32;
	qsin_lut[4805] =  9'sd37;
	icos_lut[4805] =  9'sd25;
	qsin_lut[4806] =  9'sd42;
	icos_lut[4806] =  9'sd17;
	qsin_lut[4807] =  9'sd44;
	icos_lut[4807] =  9'sd9;
	qsin_lut[4808] =  9'sd45;
	icos_lut[4808] =  9'sd0;
	qsin_lut[4809] =  9'sd44;
	icos_lut[4809] = -9'sd9;
	qsin_lut[4810] =  9'sd42;
	icos_lut[4810] = -9'sd17;
	qsin_lut[4811] =  9'sd37;
	icos_lut[4811] = -9'sd25;
	qsin_lut[4812] =  9'sd32;
	icos_lut[4812] = -9'sd32;
	qsin_lut[4813] =  9'sd25;
	icos_lut[4813] = -9'sd37;
	qsin_lut[4814] =  9'sd17;
	icos_lut[4814] = -9'sd42;
	qsin_lut[4815] =  9'sd9;
	icos_lut[4815] = -9'sd44;
	qsin_lut[4816] =  9'sd0;
	icos_lut[4816] = -9'sd45;
	qsin_lut[4817] = -9'sd9;
	icos_lut[4817] = -9'sd44;
	qsin_lut[4818] = -9'sd17;
	icos_lut[4818] = -9'sd42;
	qsin_lut[4819] = -9'sd25;
	icos_lut[4819] = -9'sd37;
	qsin_lut[4820] = -9'sd32;
	icos_lut[4820] = -9'sd32;
	qsin_lut[4821] = -9'sd37;
	icos_lut[4821] = -9'sd25;
	qsin_lut[4822] = -9'sd42;
	icos_lut[4822] = -9'sd17;
	qsin_lut[4823] = -9'sd44;
	icos_lut[4823] = -9'sd9;
	qsin_lut[4824] = -9'sd45;
	icos_lut[4824] = -9'sd0;
	qsin_lut[4825] = -9'sd44;
	icos_lut[4825] =  9'sd9;
	qsin_lut[4826] = -9'sd42;
	icos_lut[4826] =  9'sd17;
	qsin_lut[4827] = -9'sd37;
	icos_lut[4827] =  9'sd25;
	qsin_lut[4828] = -9'sd32;
	icos_lut[4828] =  9'sd32;
	qsin_lut[4829] = -9'sd25;
	icos_lut[4829] =  9'sd37;
	qsin_lut[4830] = -9'sd17;
	icos_lut[4830] =  9'sd42;
	qsin_lut[4831] = -9'sd9;
	icos_lut[4831] =  9'sd44;
	qsin_lut[4832] =  9'sd0;
	icos_lut[4832] =  9'sd47;
	qsin_lut[4833] =  9'sd9;
	icos_lut[4833] =  9'sd46;
	qsin_lut[4834] =  9'sd18;
	icos_lut[4834] =  9'sd43;
	qsin_lut[4835] =  9'sd26;
	icos_lut[4835] =  9'sd39;
	qsin_lut[4836] =  9'sd33;
	icos_lut[4836] =  9'sd33;
	qsin_lut[4837] =  9'sd39;
	icos_lut[4837] =  9'sd26;
	qsin_lut[4838] =  9'sd43;
	icos_lut[4838] =  9'sd18;
	qsin_lut[4839] =  9'sd46;
	icos_lut[4839] =  9'sd9;
	qsin_lut[4840] =  9'sd47;
	icos_lut[4840] =  9'sd0;
	qsin_lut[4841] =  9'sd46;
	icos_lut[4841] = -9'sd9;
	qsin_lut[4842] =  9'sd43;
	icos_lut[4842] = -9'sd18;
	qsin_lut[4843] =  9'sd39;
	icos_lut[4843] = -9'sd26;
	qsin_lut[4844] =  9'sd33;
	icos_lut[4844] = -9'sd33;
	qsin_lut[4845] =  9'sd26;
	icos_lut[4845] = -9'sd39;
	qsin_lut[4846] =  9'sd18;
	icos_lut[4846] = -9'sd43;
	qsin_lut[4847] =  9'sd9;
	icos_lut[4847] = -9'sd46;
	qsin_lut[4848] =  9'sd0;
	icos_lut[4848] = -9'sd47;
	qsin_lut[4849] = -9'sd9;
	icos_lut[4849] = -9'sd46;
	qsin_lut[4850] = -9'sd18;
	icos_lut[4850] = -9'sd43;
	qsin_lut[4851] = -9'sd26;
	icos_lut[4851] = -9'sd39;
	qsin_lut[4852] = -9'sd33;
	icos_lut[4852] = -9'sd33;
	qsin_lut[4853] = -9'sd39;
	icos_lut[4853] = -9'sd26;
	qsin_lut[4854] = -9'sd43;
	icos_lut[4854] = -9'sd18;
	qsin_lut[4855] = -9'sd46;
	icos_lut[4855] = -9'sd9;
	qsin_lut[4856] = -9'sd47;
	icos_lut[4856] = -9'sd0;
	qsin_lut[4857] = -9'sd46;
	icos_lut[4857] =  9'sd9;
	qsin_lut[4858] = -9'sd43;
	icos_lut[4858] =  9'sd18;
	qsin_lut[4859] = -9'sd39;
	icos_lut[4859] =  9'sd26;
	qsin_lut[4860] = -9'sd33;
	icos_lut[4860] =  9'sd33;
	qsin_lut[4861] = -9'sd26;
	icos_lut[4861] =  9'sd39;
	qsin_lut[4862] = -9'sd18;
	icos_lut[4862] =  9'sd43;
	qsin_lut[4863] = -9'sd9;
	icos_lut[4863] =  9'sd46;
	qsin_lut[4864] =  9'sd0;
	icos_lut[4864] =  9'sd49;
	qsin_lut[4865] =  9'sd10;
	icos_lut[4865] =  9'sd48;
	qsin_lut[4866] =  9'sd19;
	icos_lut[4866] =  9'sd45;
	qsin_lut[4867] =  9'sd27;
	icos_lut[4867] =  9'sd41;
	qsin_lut[4868] =  9'sd35;
	icos_lut[4868] =  9'sd35;
	qsin_lut[4869] =  9'sd41;
	icos_lut[4869] =  9'sd27;
	qsin_lut[4870] =  9'sd45;
	icos_lut[4870] =  9'sd19;
	qsin_lut[4871] =  9'sd48;
	icos_lut[4871] =  9'sd10;
	qsin_lut[4872] =  9'sd49;
	icos_lut[4872] =  9'sd0;
	qsin_lut[4873] =  9'sd48;
	icos_lut[4873] = -9'sd10;
	qsin_lut[4874] =  9'sd45;
	icos_lut[4874] = -9'sd19;
	qsin_lut[4875] =  9'sd41;
	icos_lut[4875] = -9'sd27;
	qsin_lut[4876] =  9'sd35;
	icos_lut[4876] = -9'sd35;
	qsin_lut[4877] =  9'sd27;
	icos_lut[4877] = -9'sd41;
	qsin_lut[4878] =  9'sd19;
	icos_lut[4878] = -9'sd45;
	qsin_lut[4879] =  9'sd10;
	icos_lut[4879] = -9'sd48;
	qsin_lut[4880] =  9'sd0;
	icos_lut[4880] = -9'sd49;
	qsin_lut[4881] = -9'sd10;
	icos_lut[4881] = -9'sd48;
	qsin_lut[4882] = -9'sd19;
	icos_lut[4882] = -9'sd45;
	qsin_lut[4883] = -9'sd27;
	icos_lut[4883] = -9'sd41;
	qsin_lut[4884] = -9'sd35;
	icos_lut[4884] = -9'sd35;
	qsin_lut[4885] = -9'sd41;
	icos_lut[4885] = -9'sd27;
	qsin_lut[4886] = -9'sd45;
	icos_lut[4886] = -9'sd19;
	qsin_lut[4887] = -9'sd48;
	icos_lut[4887] = -9'sd10;
	qsin_lut[4888] = -9'sd49;
	icos_lut[4888] = -9'sd0;
	qsin_lut[4889] = -9'sd48;
	icos_lut[4889] =  9'sd10;
	qsin_lut[4890] = -9'sd45;
	icos_lut[4890] =  9'sd19;
	qsin_lut[4891] = -9'sd41;
	icos_lut[4891] =  9'sd27;
	qsin_lut[4892] = -9'sd35;
	icos_lut[4892] =  9'sd35;
	qsin_lut[4893] = -9'sd27;
	icos_lut[4893] =  9'sd41;
	qsin_lut[4894] = -9'sd19;
	icos_lut[4894] =  9'sd45;
	qsin_lut[4895] = -9'sd10;
	icos_lut[4895] =  9'sd48;
	qsin_lut[4896] =  9'sd0;
	icos_lut[4896] =  9'sd51;
	qsin_lut[4897] =  9'sd10;
	icos_lut[4897] =  9'sd50;
	qsin_lut[4898] =  9'sd20;
	icos_lut[4898] =  9'sd47;
	qsin_lut[4899] =  9'sd28;
	icos_lut[4899] =  9'sd42;
	qsin_lut[4900] =  9'sd36;
	icos_lut[4900] =  9'sd36;
	qsin_lut[4901] =  9'sd42;
	icos_lut[4901] =  9'sd28;
	qsin_lut[4902] =  9'sd47;
	icos_lut[4902] =  9'sd20;
	qsin_lut[4903] =  9'sd50;
	icos_lut[4903] =  9'sd10;
	qsin_lut[4904] =  9'sd51;
	icos_lut[4904] =  9'sd0;
	qsin_lut[4905] =  9'sd50;
	icos_lut[4905] = -9'sd10;
	qsin_lut[4906] =  9'sd47;
	icos_lut[4906] = -9'sd20;
	qsin_lut[4907] =  9'sd42;
	icos_lut[4907] = -9'sd28;
	qsin_lut[4908] =  9'sd36;
	icos_lut[4908] = -9'sd36;
	qsin_lut[4909] =  9'sd28;
	icos_lut[4909] = -9'sd42;
	qsin_lut[4910] =  9'sd20;
	icos_lut[4910] = -9'sd47;
	qsin_lut[4911] =  9'sd10;
	icos_lut[4911] = -9'sd50;
	qsin_lut[4912] =  9'sd0;
	icos_lut[4912] = -9'sd51;
	qsin_lut[4913] = -9'sd10;
	icos_lut[4913] = -9'sd50;
	qsin_lut[4914] = -9'sd20;
	icos_lut[4914] = -9'sd47;
	qsin_lut[4915] = -9'sd28;
	icos_lut[4915] = -9'sd42;
	qsin_lut[4916] = -9'sd36;
	icos_lut[4916] = -9'sd36;
	qsin_lut[4917] = -9'sd42;
	icos_lut[4917] = -9'sd28;
	qsin_lut[4918] = -9'sd47;
	icos_lut[4918] = -9'sd20;
	qsin_lut[4919] = -9'sd50;
	icos_lut[4919] = -9'sd10;
	qsin_lut[4920] = -9'sd51;
	icos_lut[4920] = -9'sd0;
	qsin_lut[4921] = -9'sd50;
	icos_lut[4921] =  9'sd10;
	qsin_lut[4922] = -9'sd47;
	icos_lut[4922] =  9'sd20;
	qsin_lut[4923] = -9'sd42;
	icos_lut[4923] =  9'sd28;
	qsin_lut[4924] = -9'sd36;
	icos_lut[4924] =  9'sd36;
	qsin_lut[4925] = -9'sd28;
	icos_lut[4925] =  9'sd42;
	qsin_lut[4926] = -9'sd20;
	icos_lut[4926] =  9'sd47;
	qsin_lut[4927] = -9'sd10;
	icos_lut[4927] =  9'sd50;
	qsin_lut[4928] =  9'sd0;
	icos_lut[4928] =  9'sd53;
	qsin_lut[4929] =  9'sd10;
	icos_lut[4929] =  9'sd52;
	qsin_lut[4930] =  9'sd20;
	icos_lut[4930] =  9'sd49;
	qsin_lut[4931] =  9'sd29;
	icos_lut[4931] =  9'sd44;
	qsin_lut[4932] =  9'sd37;
	icos_lut[4932] =  9'sd37;
	qsin_lut[4933] =  9'sd44;
	icos_lut[4933] =  9'sd29;
	qsin_lut[4934] =  9'sd49;
	icos_lut[4934] =  9'sd20;
	qsin_lut[4935] =  9'sd52;
	icos_lut[4935] =  9'sd10;
	qsin_lut[4936] =  9'sd53;
	icos_lut[4936] =  9'sd0;
	qsin_lut[4937] =  9'sd52;
	icos_lut[4937] = -9'sd10;
	qsin_lut[4938] =  9'sd49;
	icos_lut[4938] = -9'sd20;
	qsin_lut[4939] =  9'sd44;
	icos_lut[4939] = -9'sd29;
	qsin_lut[4940] =  9'sd37;
	icos_lut[4940] = -9'sd37;
	qsin_lut[4941] =  9'sd29;
	icos_lut[4941] = -9'sd44;
	qsin_lut[4942] =  9'sd20;
	icos_lut[4942] = -9'sd49;
	qsin_lut[4943] =  9'sd10;
	icos_lut[4943] = -9'sd52;
	qsin_lut[4944] =  9'sd0;
	icos_lut[4944] = -9'sd53;
	qsin_lut[4945] = -9'sd10;
	icos_lut[4945] = -9'sd52;
	qsin_lut[4946] = -9'sd20;
	icos_lut[4946] = -9'sd49;
	qsin_lut[4947] = -9'sd29;
	icos_lut[4947] = -9'sd44;
	qsin_lut[4948] = -9'sd37;
	icos_lut[4948] = -9'sd37;
	qsin_lut[4949] = -9'sd44;
	icos_lut[4949] = -9'sd29;
	qsin_lut[4950] = -9'sd49;
	icos_lut[4950] = -9'sd20;
	qsin_lut[4951] = -9'sd52;
	icos_lut[4951] = -9'sd10;
	qsin_lut[4952] = -9'sd53;
	icos_lut[4952] = -9'sd0;
	qsin_lut[4953] = -9'sd52;
	icos_lut[4953] =  9'sd10;
	qsin_lut[4954] = -9'sd49;
	icos_lut[4954] =  9'sd20;
	qsin_lut[4955] = -9'sd44;
	icos_lut[4955] =  9'sd29;
	qsin_lut[4956] = -9'sd37;
	icos_lut[4956] =  9'sd37;
	qsin_lut[4957] = -9'sd29;
	icos_lut[4957] =  9'sd44;
	qsin_lut[4958] = -9'sd20;
	icos_lut[4958] =  9'sd49;
	qsin_lut[4959] = -9'sd10;
	icos_lut[4959] =  9'sd52;
	qsin_lut[4960] =  9'sd0;
	icos_lut[4960] =  9'sd55;
	qsin_lut[4961] =  9'sd11;
	icos_lut[4961] =  9'sd54;
	qsin_lut[4962] =  9'sd21;
	icos_lut[4962] =  9'sd51;
	qsin_lut[4963] =  9'sd31;
	icos_lut[4963] =  9'sd46;
	qsin_lut[4964] =  9'sd39;
	icos_lut[4964] =  9'sd39;
	qsin_lut[4965] =  9'sd46;
	icos_lut[4965] =  9'sd31;
	qsin_lut[4966] =  9'sd51;
	icos_lut[4966] =  9'sd21;
	qsin_lut[4967] =  9'sd54;
	icos_lut[4967] =  9'sd11;
	qsin_lut[4968] =  9'sd55;
	icos_lut[4968] =  9'sd0;
	qsin_lut[4969] =  9'sd54;
	icos_lut[4969] = -9'sd11;
	qsin_lut[4970] =  9'sd51;
	icos_lut[4970] = -9'sd21;
	qsin_lut[4971] =  9'sd46;
	icos_lut[4971] = -9'sd31;
	qsin_lut[4972] =  9'sd39;
	icos_lut[4972] = -9'sd39;
	qsin_lut[4973] =  9'sd31;
	icos_lut[4973] = -9'sd46;
	qsin_lut[4974] =  9'sd21;
	icos_lut[4974] = -9'sd51;
	qsin_lut[4975] =  9'sd11;
	icos_lut[4975] = -9'sd54;
	qsin_lut[4976] =  9'sd0;
	icos_lut[4976] = -9'sd55;
	qsin_lut[4977] = -9'sd11;
	icos_lut[4977] = -9'sd54;
	qsin_lut[4978] = -9'sd21;
	icos_lut[4978] = -9'sd51;
	qsin_lut[4979] = -9'sd31;
	icos_lut[4979] = -9'sd46;
	qsin_lut[4980] = -9'sd39;
	icos_lut[4980] = -9'sd39;
	qsin_lut[4981] = -9'sd46;
	icos_lut[4981] = -9'sd31;
	qsin_lut[4982] = -9'sd51;
	icos_lut[4982] = -9'sd21;
	qsin_lut[4983] = -9'sd54;
	icos_lut[4983] = -9'sd11;
	qsin_lut[4984] = -9'sd55;
	icos_lut[4984] = -9'sd0;
	qsin_lut[4985] = -9'sd54;
	icos_lut[4985] =  9'sd11;
	qsin_lut[4986] = -9'sd51;
	icos_lut[4986] =  9'sd21;
	qsin_lut[4987] = -9'sd46;
	icos_lut[4987] =  9'sd31;
	qsin_lut[4988] = -9'sd39;
	icos_lut[4988] =  9'sd39;
	qsin_lut[4989] = -9'sd31;
	icos_lut[4989] =  9'sd46;
	qsin_lut[4990] = -9'sd21;
	icos_lut[4990] =  9'sd51;
	qsin_lut[4991] = -9'sd11;
	icos_lut[4991] =  9'sd54;
	qsin_lut[4992] =  9'sd0;
	icos_lut[4992] =  9'sd57;
	qsin_lut[4993] =  9'sd11;
	icos_lut[4993] =  9'sd56;
	qsin_lut[4994] =  9'sd22;
	icos_lut[4994] =  9'sd53;
	qsin_lut[4995] =  9'sd32;
	icos_lut[4995] =  9'sd47;
	qsin_lut[4996] =  9'sd40;
	icos_lut[4996] =  9'sd40;
	qsin_lut[4997] =  9'sd47;
	icos_lut[4997] =  9'sd32;
	qsin_lut[4998] =  9'sd53;
	icos_lut[4998] =  9'sd22;
	qsin_lut[4999] =  9'sd56;
	icos_lut[4999] =  9'sd11;
	qsin_lut[5000] =  9'sd57;
	icos_lut[5000] =  9'sd0;
	qsin_lut[5001] =  9'sd56;
	icos_lut[5001] = -9'sd11;
	qsin_lut[5002] =  9'sd53;
	icos_lut[5002] = -9'sd22;
	qsin_lut[5003] =  9'sd47;
	icos_lut[5003] = -9'sd32;
	qsin_lut[5004] =  9'sd40;
	icos_lut[5004] = -9'sd40;
	qsin_lut[5005] =  9'sd32;
	icos_lut[5005] = -9'sd47;
	qsin_lut[5006] =  9'sd22;
	icos_lut[5006] = -9'sd53;
	qsin_lut[5007] =  9'sd11;
	icos_lut[5007] = -9'sd56;
	qsin_lut[5008] =  9'sd0;
	icos_lut[5008] = -9'sd57;
	qsin_lut[5009] = -9'sd11;
	icos_lut[5009] = -9'sd56;
	qsin_lut[5010] = -9'sd22;
	icos_lut[5010] = -9'sd53;
	qsin_lut[5011] = -9'sd32;
	icos_lut[5011] = -9'sd47;
	qsin_lut[5012] = -9'sd40;
	icos_lut[5012] = -9'sd40;
	qsin_lut[5013] = -9'sd47;
	icos_lut[5013] = -9'sd32;
	qsin_lut[5014] = -9'sd53;
	icos_lut[5014] = -9'sd22;
	qsin_lut[5015] = -9'sd56;
	icos_lut[5015] = -9'sd11;
	qsin_lut[5016] = -9'sd57;
	icos_lut[5016] = -9'sd0;
	qsin_lut[5017] = -9'sd56;
	icos_lut[5017] =  9'sd11;
	qsin_lut[5018] = -9'sd53;
	icos_lut[5018] =  9'sd22;
	qsin_lut[5019] = -9'sd47;
	icos_lut[5019] =  9'sd32;
	qsin_lut[5020] = -9'sd40;
	icos_lut[5020] =  9'sd40;
	qsin_lut[5021] = -9'sd32;
	icos_lut[5021] =  9'sd47;
	qsin_lut[5022] = -9'sd22;
	icos_lut[5022] =  9'sd53;
	qsin_lut[5023] = -9'sd11;
	icos_lut[5023] =  9'sd56;
	qsin_lut[5024] =  9'sd0;
	icos_lut[5024] =  9'sd59;
	qsin_lut[5025] =  9'sd12;
	icos_lut[5025] =  9'sd58;
	qsin_lut[5026] =  9'sd23;
	icos_lut[5026] =  9'sd55;
	qsin_lut[5027] =  9'sd33;
	icos_lut[5027] =  9'sd49;
	qsin_lut[5028] =  9'sd42;
	icos_lut[5028] =  9'sd42;
	qsin_lut[5029] =  9'sd49;
	icos_lut[5029] =  9'sd33;
	qsin_lut[5030] =  9'sd55;
	icos_lut[5030] =  9'sd23;
	qsin_lut[5031] =  9'sd58;
	icos_lut[5031] =  9'sd12;
	qsin_lut[5032] =  9'sd59;
	icos_lut[5032] =  9'sd0;
	qsin_lut[5033] =  9'sd58;
	icos_lut[5033] = -9'sd12;
	qsin_lut[5034] =  9'sd55;
	icos_lut[5034] = -9'sd23;
	qsin_lut[5035] =  9'sd49;
	icos_lut[5035] = -9'sd33;
	qsin_lut[5036] =  9'sd42;
	icos_lut[5036] = -9'sd42;
	qsin_lut[5037] =  9'sd33;
	icos_lut[5037] = -9'sd49;
	qsin_lut[5038] =  9'sd23;
	icos_lut[5038] = -9'sd55;
	qsin_lut[5039] =  9'sd12;
	icos_lut[5039] = -9'sd58;
	qsin_lut[5040] =  9'sd0;
	icos_lut[5040] = -9'sd59;
	qsin_lut[5041] = -9'sd12;
	icos_lut[5041] = -9'sd58;
	qsin_lut[5042] = -9'sd23;
	icos_lut[5042] = -9'sd55;
	qsin_lut[5043] = -9'sd33;
	icos_lut[5043] = -9'sd49;
	qsin_lut[5044] = -9'sd42;
	icos_lut[5044] = -9'sd42;
	qsin_lut[5045] = -9'sd49;
	icos_lut[5045] = -9'sd33;
	qsin_lut[5046] = -9'sd55;
	icos_lut[5046] = -9'sd23;
	qsin_lut[5047] = -9'sd58;
	icos_lut[5047] = -9'sd12;
	qsin_lut[5048] = -9'sd59;
	icos_lut[5048] = -9'sd0;
	qsin_lut[5049] = -9'sd58;
	icos_lut[5049] =  9'sd12;
	qsin_lut[5050] = -9'sd55;
	icos_lut[5050] =  9'sd23;
	qsin_lut[5051] = -9'sd49;
	icos_lut[5051] =  9'sd33;
	qsin_lut[5052] = -9'sd42;
	icos_lut[5052] =  9'sd42;
	qsin_lut[5053] = -9'sd33;
	icos_lut[5053] =  9'sd49;
	qsin_lut[5054] = -9'sd23;
	icos_lut[5054] =  9'sd55;
	qsin_lut[5055] = -9'sd12;
	icos_lut[5055] =  9'sd58;
	qsin_lut[5056] =  9'sd0;
	icos_lut[5056] =  9'sd61;
	qsin_lut[5057] =  9'sd12;
	icos_lut[5057] =  9'sd60;
	qsin_lut[5058] =  9'sd23;
	icos_lut[5058] =  9'sd56;
	qsin_lut[5059] =  9'sd34;
	icos_lut[5059] =  9'sd51;
	qsin_lut[5060] =  9'sd43;
	icos_lut[5060] =  9'sd43;
	qsin_lut[5061] =  9'sd51;
	icos_lut[5061] =  9'sd34;
	qsin_lut[5062] =  9'sd56;
	icos_lut[5062] =  9'sd23;
	qsin_lut[5063] =  9'sd60;
	icos_lut[5063] =  9'sd12;
	qsin_lut[5064] =  9'sd61;
	icos_lut[5064] =  9'sd0;
	qsin_lut[5065] =  9'sd60;
	icos_lut[5065] = -9'sd12;
	qsin_lut[5066] =  9'sd56;
	icos_lut[5066] = -9'sd23;
	qsin_lut[5067] =  9'sd51;
	icos_lut[5067] = -9'sd34;
	qsin_lut[5068] =  9'sd43;
	icos_lut[5068] = -9'sd43;
	qsin_lut[5069] =  9'sd34;
	icos_lut[5069] = -9'sd51;
	qsin_lut[5070] =  9'sd23;
	icos_lut[5070] = -9'sd56;
	qsin_lut[5071] =  9'sd12;
	icos_lut[5071] = -9'sd60;
	qsin_lut[5072] =  9'sd0;
	icos_lut[5072] = -9'sd61;
	qsin_lut[5073] = -9'sd12;
	icos_lut[5073] = -9'sd60;
	qsin_lut[5074] = -9'sd23;
	icos_lut[5074] = -9'sd56;
	qsin_lut[5075] = -9'sd34;
	icos_lut[5075] = -9'sd51;
	qsin_lut[5076] = -9'sd43;
	icos_lut[5076] = -9'sd43;
	qsin_lut[5077] = -9'sd51;
	icos_lut[5077] = -9'sd34;
	qsin_lut[5078] = -9'sd56;
	icos_lut[5078] = -9'sd23;
	qsin_lut[5079] = -9'sd60;
	icos_lut[5079] = -9'sd12;
	qsin_lut[5080] = -9'sd61;
	icos_lut[5080] = -9'sd0;
	qsin_lut[5081] = -9'sd60;
	icos_lut[5081] =  9'sd12;
	qsin_lut[5082] = -9'sd56;
	icos_lut[5082] =  9'sd23;
	qsin_lut[5083] = -9'sd51;
	icos_lut[5083] =  9'sd34;
	qsin_lut[5084] = -9'sd43;
	icos_lut[5084] =  9'sd43;
	qsin_lut[5085] = -9'sd34;
	icos_lut[5085] =  9'sd51;
	qsin_lut[5086] = -9'sd23;
	icos_lut[5086] =  9'sd56;
	qsin_lut[5087] = -9'sd12;
	icos_lut[5087] =  9'sd60;
	qsin_lut[5088] =  9'sd0;
	icos_lut[5088] =  9'sd63;
	qsin_lut[5089] =  9'sd12;
	icos_lut[5089] =  9'sd62;
	qsin_lut[5090] =  9'sd24;
	icos_lut[5090] =  9'sd58;
	qsin_lut[5091] =  9'sd35;
	icos_lut[5091] =  9'sd52;
	qsin_lut[5092] =  9'sd45;
	icos_lut[5092] =  9'sd45;
	qsin_lut[5093] =  9'sd52;
	icos_lut[5093] =  9'sd35;
	qsin_lut[5094] =  9'sd58;
	icos_lut[5094] =  9'sd24;
	qsin_lut[5095] =  9'sd62;
	icos_lut[5095] =  9'sd12;
	qsin_lut[5096] =  9'sd63;
	icos_lut[5096] =  9'sd0;
	qsin_lut[5097] =  9'sd62;
	icos_lut[5097] = -9'sd12;
	qsin_lut[5098] =  9'sd58;
	icos_lut[5098] = -9'sd24;
	qsin_lut[5099] =  9'sd52;
	icos_lut[5099] = -9'sd35;
	qsin_lut[5100] =  9'sd45;
	icos_lut[5100] = -9'sd45;
	qsin_lut[5101] =  9'sd35;
	icos_lut[5101] = -9'sd52;
	qsin_lut[5102] =  9'sd24;
	icos_lut[5102] = -9'sd58;
	qsin_lut[5103] =  9'sd12;
	icos_lut[5103] = -9'sd62;
	qsin_lut[5104] =  9'sd0;
	icos_lut[5104] = -9'sd63;
	qsin_lut[5105] = -9'sd12;
	icos_lut[5105] = -9'sd62;
	qsin_lut[5106] = -9'sd24;
	icos_lut[5106] = -9'sd58;
	qsin_lut[5107] = -9'sd35;
	icos_lut[5107] = -9'sd52;
	qsin_lut[5108] = -9'sd45;
	icos_lut[5108] = -9'sd45;
	qsin_lut[5109] = -9'sd52;
	icos_lut[5109] = -9'sd35;
	qsin_lut[5110] = -9'sd58;
	icos_lut[5110] = -9'sd24;
	qsin_lut[5111] = -9'sd62;
	icos_lut[5111] = -9'sd12;
	qsin_lut[5112] = -9'sd63;
	icos_lut[5112] = -9'sd0;
	qsin_lut[5113] = -9'sd62;
	icos_lut[5113] =  9'sd12;
	qsin_lut[5114] = -9'sd58;
	icos_lut[5114] =  9'sd24;
	qsin_lut[5115] = -9'sd52;
	icos_lut[5115] =  9'sd35;
	qsin_lut[5116] = -9'sd45;
	icos_lut[5116] =  9'sd45;
	qsin_lut[5117] = -9'sd35;
	icos_lut[5117] =  9'sd52;
	qsin_lut[5118] = -9'sd24;
	icos_lut[5118] =  9'sd58;
	qsin_lut[5119] = -9'sd12;
	icos_lut[5119] =  9'sd62;
	qsin_lut[5120] =  9'sd0;
	icos_lut[5120] =  9'sd65;
	qsin_lut[5121] =  9'sd13;
	icos_lut[5121] =  9'sd64;
	qsin_lut[5122] =  9'sd25;
	icos_lut[5122] =  9'sd60;
	qsin_lut[5123] =  9'sd36;
	icos_lut[5123] =  9'sd54;
	qsin_lut[5124] =  9'sd46;
	icos_lut[5124] =  9'sd46;
	qsin_lut[5125] =  9'sd54;
	icos_lut[5125] =  9'sd36;
	qsin_lut[5126] =  9'sd60;
	icos_lut[5126] =  9'sd25;
	qsin_lut[5127] =  9'sd64;
	icos_lut[5127] =  9'sd13;
	qsin_lut[5128] =  9'sd65;
	icos_lut[5128] =  9'sd0;
	qsin_lut[5129] =  9'sd64;
	icos_lut[5129] = -9'sd13;
	qsin_lut[5130] =  9'sd60;
	icos_lut[5130] = -9'sd25;
	qsin_lut[5131] =  9'sd54;
	icos_lut[5131] = -9'sd36;
	qsin_lut[5132] =  9'sd46;
	icos_lut[5132] = -9'sd46;
	qsin_lut[5133] =  9'sd36;
	icos_lut[5133] = -9'sd54;
	qsin_lut[5134] =  9'sd25;
	icos_lut[5134] = -9'sd60;
	qsin_lut[5135] =  9'sd13;
	icos_lut[5135] = -9'sd64;
	qsin_lut[5136] =  9'sd0;
	icos_lut[5136] = -9'sd65;
	qsin_lut[5137] = -9'sd13;
	icos_lut[5137] = -9'sd64;
	qsin_lut[5138] = -9'sd25;
	icos_lut[5138] = -9'sd60;
	qsin_lut[5139] = -9'sd36;
	icos_lut[5139] = -9'sd54;
	qsin_lut[5140] = -9'sd46;
	icos_lut[5140] = -9'sd46;
	qsin_lut[5141] = -9'sd54;
	icos_lut[5141] = -9'sd36;
	qsin_lut[5142] = -9'sd60;
	icos_lut[5142] = -9'sd25;
	qsin_lut[5143] = -9'sd64;
	icos_lut[5143] = -9'sd13;
	qsin_lut[5144] = -9'sd65;
	icos_lut[5144] = -9'sd0;
	qsin_lut[5145] = -9'sd64;
	icos_lut[5145] =  9'sd13;
	qsin_lut[5146] = -9'sd60;
	icos_lut[5146] =  9'sd25;
	qsin_lut[5147] = -9'sd54;
	icos_lut[5147] =  9'sd36;
	qsin_lut[5148] = -9'sd46;
	icos_lut[5148] =  9'sd46;
	qsin_lut[5149] = -9'sd36;
	icos_lut[5149] =  9'sd54;
	qsin_lut[5150] = -9'sd25;
	icos_lut[5150] =  9'sd60;
	qsin_lut[5151] = -9'sd13;
	icos_lut[5151] =  9'sd64;
	qsin_lut[5152] =  9'sd0;
	icos_lut[5152] =  9'sd67;
	qsin_lut[5153] =  9'sd13;
	icos_lut[5153] =  9'sd66;
	qsin_lut[5154] =  9'sd26;
	icos_lut[5154] =  9'sd62;
	qsin_lut[5155] =  9'sd37;
	icos_lut[5155] =  9'sd56;
	qsin_lut[5156] =  9'sd47;
	icos_lut[5156] =  9'sd47;
	qsin_lut[5157] =  9'sd56;
	icos_lut[5157] =  9'sd37;
	qsin_lut[5158] =  9'sd62;
	icos_lut[5158] =  9'sd26;
	qsin_lut[5159] =  9'sd66;
	icos_lut[5159] =  9'sd13;
	qsin_lut[5160] =  9'sd67;
	icos_lut[5160] =  9'sd0;
	qsin_lut[5161] =  9'sd66;
	icos_lut[5161] = -9'sd13;
	qsin_lut[5162] =  9'sd62;
	icos_lut[5162] = -9'sd26;
	qsin_lut[5163] =  9'sd56;
	icos_lut[5163] = -9'sd37;
	qsin_lut[5164] =  9'sd47;
	icos_lut[5164] = -9'sd47;
	qsin_lut[5165] =  9'sd37;
	icos_lut[5165] = -9'sd56;
	qsin_lut[5166] =  9'sd26;
	icos_lut[5166] = -9'sd62;
	qsin_lut[5167] =  9'sd13;
	icos_lut[5167] = -9'sd66;
	qsin_lut[5168] =  9'sd0;
	icos_lut[5168] = -9'sd67;
	qsin_lut[5169] = -9'sd13;
	icos_lut[5169] = -9'sd66;
	qsin_lut[5170] = -9'sd26;
	icos_lut[5170] = -9'sd62;
	qsin_lut[5171] = -9'sd37;
	icos_lut[5171] = -9'sd56;
	qsin_lut[5172] = -9'sd47;
	icos_lut[5172] = -9'sd47;
	qsin_lut[5173] = -9'sd56;
	icos_lut[5173] = -9'sd37;
	qsin_lut[5174] = -9'sd62;
	icos_lut[5174] = -9'sd26;
	qsin_lut[5175] = -9'sd66;
	icos_lut[5175] = -9'sd13;
	qsin_lut[5176] = -9'sd67;
	icos_lut[5176] = -9'sd0;
	qsin_lut[5177] = -9'sd66;
	icos_lut[5177] =  9'sd13;
	qsin_lut[5178] = -9'sd62;
	icos_lut[5178] =  9'sd26;
	qsin_lut[5179] = -9'sd56;
	icos_lut[5179] =  9'sd37;
	qsin_lut[5180] = -9'sd47;
	icos_lut[5180] =  9'sd47;
	qsin_lut[5181] = -9'sd37;
	icos_lut[5181] =  9'sd56;
	qsin_lut[5182] = -9'sd26;
	icos_lut[5182] =  9'sd62;
	qsin_lut[5183] = -9'sd13;
	icos_lut[5183] =  9'sd66;
	qsin_lut[5184] =  9'sd0;
	icos_lut[5184] =  9'sd69;
	qsin_lut[5185] =  9'sd13;
	icos_lut[5185] =  9'sd68;
	qsin_lut[5186] =  9'sd26;
	icos_lut[5186] =  9'sd64;
	qsin_lut[5187] =  9'sd38;
	icos_lut[5187] =  9'sd57;
	qsin_lut[5188] =  9'sd49;
	icos_lut[5188] =  9'sd49;
	qsin_lut[5189] =  9'sd57;
	icos_lut[5189] =  9'sd38;
	qsin_lut[5190] =  9'sd64;
	icos_lut[5190] =  9'sd26;
	qsin_lut[5191] =  9'sd68;
	icos_lut[5191] =  9'sd13;
	qsin_lut[5192] =  9'sd69;
	icos_lut[5192] =  9'sd0;
	qsin_lut[5193] =  9'sd68;
	icos_lut[5193] = -9'sd13;
	qsin_lut[5194] =  9'sd64;
	icos_lut[5194] = -9'sd26;
	qsin_lut[5195] =  9'sd57;
	icos_lut[5195] = -9'sd38;
	qsin_lut[5196] =  9'sd49;
	icos_lut[5196] = -9'sd49;
	qsin_lut[5197] =  9'sd38;
	icos_lut[5197] = -9'sd57;
	qsin_lut[5198] =  9'sd26;
	icos_lut[5198] = -9'sd64;
	qsin_lut[5199] =  9'sd13;
	icos_lut[5199] = -9'sd68;
	qsin_lut[5200] =  9'sd0;
	icos_lut[5200] = -9'sd69;
	qsin_lut[5201] = -9'sd13;
	icos_lut[5201] = -9'sd68;
	qsin_lut[5202] = -9'sd26;
	icos_lut[5202] = -9'sd64;
	qsin_lut[5203] = -9'sd38;
	icos_lut[5203] = -9'sd57;
	qsin_lut[5204] = -9'sd49;
	icos_lut[5204] = -9'sd49;
	qsin_lut[5205] = -9'sd57;
	icos_lut[5205] = -9'sd38;
	qsin_lut[5206] = -9'sd64;
	icos_lut[5206] = -9'sd26;
	qsin_lut[5207] = -9'sd68;
	icos_lut[5207] = -9'sd13;
	qsin_lut[5208] = -9'sd69;
	icos_lut[5208] = -9'sd0;
	qsin_lut[5209] = -9'sd68;
	icos_lut[5209] =  9'sd13;
	qsin_lut[5210] = -9'sd64;
	icos_lut[5210] =  9'sd26;
	qsin_lut[5211] = -9'sd57;
	icos_lut[5211] =  9'sd38;
	qsin_lut[5212] = -9'sd49;
	icos_lut[5212] =  9'sd49;
	qsin_lut[5213] = -9'sd38;
	icos_lut[5213] =  9'sd57;
	qsin_lut[5214] = -9'sd26;
	icos_lut[5214] =  9'sd64;
	qsin_lut[5215] = -9'sd13;
	icos_lut[5215] =  9'sd68;
	qsin_lut[5216] =  9'sd0;
	icos_lut[5216] =  9'sd71;
	qsin_lut[5217] =  9'sd14;
	icos_lut[5217] =  9'sd70;
	qsin_lut[5218] =  9'sd27;
	icos_lut[5218] =  9'sd66;
	qsin_lut[5219] =  9'sd39;
	icos_lut[5219] =  9'sd59;
	qsin_lut[5220] =  9'sd50;
	icos_lut[5220] =  9'sd50;
	qsin_lut[5221] =  9'sd59;
	icos_lut[5221] =  9'sd39;
	qsin_lut[5222] =  9'sd66;
	icos_lut[5222] =  9'sd27;
	qsin_lut[5223] =  9'sd70;
	icos_lut[5223] =  9'sd14;
	qsin_lut[5224] =  9'sd71;
	icos_lut[5224] =  9'sd0;
	qsin_lut[5225] =  9'sd70;
	icos_lut[5225] = -9'sd14;
	qsin_lut[5226] =  9'sd66;
	icos_lut[5226] = -9'sd27;
	qsin_lut[5227] =  9'sd59;
	icos_lut[5227] = -9'sd39;
	qsin_lut[5228] =  9'sd50;
	icos_lut[5228] = -9'sd50;
	qsin_lut[5229] =  9'sd39;
	icos_lut[5229] = -9'sd59;
	qsin_lut[5230] =  9'sd27;
	icos_lut[5230] = -9'sd66;
	qsin_lut[5231] =  9'sd14;
	icos_lut[5231] = -9'sd70;
	qsin_lut[5232] =  9'sd0;
	icos_lut[5232] = -9'sd71;
	qsin_lut[5233] = -9'sd14;
	icos_lut[5233] = -9'sd70;
	qsin_lut[5234] = -9'sd27;
	icos_lut[5234] = -9'sd66;
	qsin_lut[5235] = -9'sd39;
	icos_lut[5235] = -9'sd59;
	qsin_lut[5236] = -9'sd50;
	icos_lut[5236] = -9'sd50;
	qsin_lut[5237] = -9'sd59;
	icos_lut[5237] = -9'sd39;
	qsin_lut[5238] = -9'sd66;
	icos_lut[5238] = -9'sd27;
	qsin_lut[5239] = -9'sd70;
	icos_lut[5239] = -9'sd14;
	qsin_lut[5240] = -9'sd71;
	icos_lut[5240] = -9'sd0;
	qsin_lut[5241] = -9'sd70;
	icos_lut[5241] =  9'sd14;
	qsin_lut[5242] = -9'sd66;
	icos_lut[5242] =  9'sd27;
	qsin_lut[5243] = -9'sd59;
	icos_lut[5243] =  9'sd39;
	qsin_lut[5244] = -9'sd50;
	icos_lut[5244] =  9'sd50;
	qsin_lut[5245] = -9'sd39;
	icos_lut[5245] =  9'sd59;
	qsin_lut[5246] = -9'sd27;
	icos_lut[5246] =  9'sd66;
	qsin_lut[5247] = -9'sd14;
	icos_lut[5247] =  9'sd70;
	qsin_lut[5248] =  9'sd0;
	icos_lut[5248] =  9'sd73;
	qsin_lut[5249] =  9'sd14;
	icos_lut[5249] =  9'sd72;
	qsin_lut[5250] =  9'sd28;
	icos_lut[5250] =  9'sd67;
	qsin_lut[5251] =  9'sd41;
	icos_lut[5251] =  9'sd61;
	qsin_lut[5252] =  9'sd52;
	icos_lut[5252] =  9'sd52;
	qsin_lut[5253] =  9'sd61;
	icos_lut[5253] =  9'sd41;
	qsin_lut[5254] =  9'sd67;
	icos_lut[5254] =  9'sd28;
	qsin_lut[5255] =  9'sd72;
	icos_lut[5255] =  9'sd14;
	qsin_lut[5256] =  9'sd73;
	icos_lut[5256] =  9'sd0;
	qsin_lut[5257] =  9'sd72;
	icos_lut[5257] = -9'sd14;
	qsin_lut[5258] =  9'sd67;
	icos_lut[5258] = -9'sd28;
	qsin_lut[5259] =  9'sd61;
	icos_lut[5259] = -9'sd41;
	qsin_lut[5260] =  9'sd52;
	icos_lut[5260] = -9'sd52;
	qsin_lut[5261] =  9'sd41;
	icos_lut[5261] = -9'sd61;
	qsin_lut[5262] =  9'sd28;
	icos_lut[5262] = -9'sd67;
	qsin_lut[5263] =  9'sd14;
	icos_lut[5263] = -9'sd72;
	qsin_lut[5264] =  9'sd0;
	icos_lut[5264] = -9'sd73;
	qsin_lut[5265] = -9'sd14;
	icos_lut[5265] = -9'sd72;
	qsin_lut[5266] = -9'sd28;
	icos_lut[5266] = -9'sd67;
	qsin_lut[5267] = -9'sd41;
	icos_lut[5267] = -9'sd61;
	qsin_lut[5268] = -9'sd52;
	icos_lut[5268] = -9'sd52;
	qsin_lut[5269] = -9'sd61;
	icos_lut[5269] = -9'sd41;
	qsin_lut[5270] = -9'sd67;
	icos_lut[5270] = -9'sd28;
	qsin_lut[5271] = -9'sd72;
	icos_lut[5271] = -9'sd14;
	qsin_lut[5272] = -9'sd73;
	icos_lut[5272] = -9'sd0;
	qsin_lut[5273] = -9'sd72;
	icos_lut[5273] =  9'sd14;
	qsin_lut[5274] = -9'sd67;
	icos_lut[5274] =  9'sd28;
	qsin_lut[5275] = -9'sd61;
	icos_lut[5275] =  9'sd41;
	qsin_lut[5276] = -9'sd52;
	icos_lut[5276] =  9'sd52;
	qsin_lut[5277] = -9'sd41;
	icos_lut[5277] =  9'sd61;
	qsin_lut[5278] = -9'sd28;
	icos_lut[5278] =  9'sd67;
	qsin_lut[5279] = -9'sd14;
	icos_lut[5279] =  9'sd72;
	qsin_lut[5280] =  9'sd0;
	icos_lut[5280] =  9'sd75;
	qsin_lut[5281] =  9'sd15;
	icos_lut[5281] =  9'sd74;
	qsin_lut[5282] =  9'sd29;
	icos_lut[5282] =  9'sd69;
	qsin_lut[5283] =  9'sd42;
	icos_lut[5283] =  9'sd62;
	qsin_lut[5284] =  9'sd53;
	icos_lut[5284] =  9'sd53;
	qsin_lut[5285] =  9'sd62;
	icos_lut[5285] =  9'sd42;
	qsin_lut[5286] =  9'sd69;
	icos_lut[5286] =  9'sd29;
	qsin_lut[5287] =  9'sd74;
	icos_lut[5287] =  9'sd15;
	qsin_lut[5288] =  9'sd75;
	icos_lut[5288] =  9'sd0;
	qsin_lut[5289] =  9'sd74;
	icos_lut[5289] = -9'sd15;
	qsin_lut[5290] =  9'sd69;
	icos_lut[5290] = -9'sd29;
	qsin_lut[5291] =  9'sd62;
	icos_lut[5291] = -9'sd42;
	qsin_lut[5292] =  9'sd53;
	icos_lut[5292] = -9'sd53;
	qsin_lut[5293] =  9'sd42;
	icos_lut[5293] = -9'sd62;
	qsin_lut[5294] =  9'sd29;
	icos_lut[5294] = -9'sd69;
	qsin_lut[5295] =  9'sd15;
	icos_lut[5295] = -9'sd74;
	qsin_lut[5296] =  9'sd0;
	icos_lut[5296] = -9'sd75;
	qsin_lut[5297] = -9'sd15;
	icos_lut[5297] = -9'sd74;
	qsin_lut[5298] = -9'sd29;
	icos_lut[5298] = -9'sd69;
	qsin_lut[5299] = -9'sd42;
	icos_lut[5299] = -9'sd62;
	qsin_lut[5300] = -9'sd53;
	icos_lut[5300] = -9'sd53;
	qsin_lut[5301] = -9'sd62;
	icos_lut[5301] = -9'sd42;
	qsin_lut[5302] = -9'sd69;
	icos_lut[5302] = -9'sd29;
	qsin_lut[5303] = -9'sd74;
	icos_lut[5303] = -9'sd15;
	qsin_lut[5304] = -9'sd75;
	icos_lut[5304] = -9'sd0;
	qsin_lut[5305] = -9'sd74;
	icos_lut[5305] =  9'sd15;
	qsin_lut[5306] = -9'sd69;
	icos_lut[5306] =  9'sd29;
	qsin_lut[5307] = -9'sd62;
	icos_lut[5307] =  9'sd42;
	qsin_lut[5308] = -9'sd53;
	icos_lut[5308] =  9'sd53;
	qsin_lut[5309] = -9'sd42;
	icos_lut[5309] =  9'sd62;
	qsin_lut[5310] = -9'sd29;
	icos_lut[5310] =  9'sd69;
	qsin_lut[5311] = -9'sd15;
	icos_lut[5311] =  9'sd74;
	qsin_lut[5312] =  9'sd0;
	icos_lut[5312] =  9'sd77;
	qsin_lut[5313] =  9'sd15;
	icos_lut[5313] =  9'sd76;
	qsin_lut[5314] =  9'sd29;
	icos_lut[5314] =  9'sd71;
	qsin_lut[5315] =  9'sd43;
	icos_lut[5315] =  9'sd64;
	qsin_lut[5316] =  9'sd54;
	icos_lut[5316] =  9'sd54;
	qsin_lut[5317] =  9'sd64;
	icos_lut[5317] =  9'sd43;
	qsin_lut[5318] =  9'sd71;
	icos_lut[5318] =  9'sd29;
	qsin_lut[5319] =  9'sd76;
	icos_lut[5319] =  9'sd15;
	qsin_lut[5320] =  9'sd77;
	icos_lut[5320] =  9'sd0;
	qsin_lut[5321] =  9'sd76;
	icos_lut[5321] = -9'sd15;
	qsin_lut[5322] =  9'sd71;
	icos_lut[5322] = -9'sd29;
	qsin_lut[5323] =  9'sd64;
	icos_lut[5323] = -9'sd43;
	qsin_lut[5324] =  9'sd54;
	icos_lut[5324] = -9'sd54;
	qsin_lut[5325] =  9'sd43;
	icos_lut[5325] = -9'sd64;
	qsin_lut[5326] =  9'sd29;
	icos_lut[5326] = -9'sd71;
	qsin_lut[5327] =  9'sd15;
	icos_lut[5327] = -9'sd76;
	qsin_lut[5328] =  9'sd0;
	icos_lut[5328] = -9'sd77;
	qsin_lut[5329] = -9'sd15;
	icos_lut[5329] = -9'sd76;
	qsin_lut[5330] = -9'sd29;
	icos_lut[5330] = -9'sd71;
	qsin_lut[5331] = -9'sd43;
	icos_lut[5331] = -9'sd64;
	qsin_lut[5332] = -9'sd54;
	icos_lut[5332] = -9'sd54;
	qsin_lut[5333] = -9'sd64;
	icos_lut[5333] = -9'sd43;
	qsin_lut[5334] = -9'sd71;
	icos_lut[5334] = -9'sd29;
	qsin_lut[5335] = -9'sd76;
	icos_lut[5335] = -9'sd15;
	qsin_lut[5336] = -9'sd77;
	icos_lut[5336] = -9'sd0;
	qsin_lut[5337] = -9'sd76;
	icos_lut[5337] =  9'sd15;
	qsin_lut[5338] = -9'sd71;
	icos_lut[5338] =  9'sd29;
	qsin_lut[5339] = -9'sd64;
	icos_lut[5339] =  9'sd43;
	qsin_lut[5340] = -9'sd54;
	icos_lut[5340] =  9'sd54;
	qsin_lut[5341] = -9'sd43;
	icos_lut[5341] =  9'sd64;
	qsin_lut[5342] = -9'sd29;
	icos_lut[5342] =  9'sd71;
	qsin_lut[5343] = -9'sd15;
	icos_lut[5343] =  9'sd76;
	qsin_lut[5344] =  9'sd0;
	icos_lut[5344] =  9'sd79;
	qsin_lut[5345] =  9'sd15;
	icos_lut[5345] =  9'sd77;
	qsin_lut[5346] =  9'sd30;
	icos_lut[5346] =  9'sd73;
	qsin_lut[5347] =  9'sd44;
	icos_lut[5347] =  9'sd66;
	qsin_lut[5348] =  9'sd56;
	icos_lut[5348] =  9'sd56;
	qsin_lut[5349] =  9'sd66;
	icos_lut[5349] =  9'sd44;
	qsin_lut[5350] =  9'sd73;
	icos_lut[5350] =  9'sd30;
	qsin_lut[5351] =  9'sd77;
	icos_lut[5351] =  9'sd15;
	qsin_lut[5352] =  9'sd79;
	icos_lut[5352] =  9'sd0;
	qsin_lut[5353] =  9'sd77;
	icos_lut[5353] = -9'sd15;
	qsin_lut[5354] =  9'sd73;
	icos_lut[5354] = -9'sd30;
	qsin_lut[5355] =  9'sd66;
	icos_lut[5355] = -9'sd44;
	qsin_lut[5356] =  9'sd56;
	icos_lut[5356] = -9'sd56;
	qsin_lut[5357] =  9'sd44;
	icos_lut[5357] = -9'sd66;
	qsin_lut[5358] =  9'sd30;
	icos_lut[5358] = -9'sd73;
	qsin_lut[5359] =  9'sd15;
	icos_lut[5359] = -9'sd77;
	qsin_lut[5360] =  9'sd0;
	icos_lut[5360] = -9'sd79;
	qsin_lut[5361] = -9'sd15;
	icos_lut[5361] = -9'sd77;
	qsin_lut[5362] = -9'sd30;
	icos_lut[5362] = -9'sd73;
	qsin_lut[5363] = -9'sd44;
	icos_lut[5363] = -9'sd66;
	qsin_lut[5364] = -9'sd56;
	icos_lut[5364] = -9'sd56;
	qsin_lut[5365] = -9'sd66;
	icos_lut[5365] = -9'sd44;
	qsin_lut[5366] = -9'sd73;
	icos_lut[5366] = -9'sd30;
	qsin_lut[5367] = -9'sd77;
	icos_lut[5367] = -9'sd15;
	qsin_lut[5368] = -9'sd79;
	icos_lut[5368] = -9'sd0;
	qsin_lut[5369] = -9'sd77;
	icos_lut[5369] =  9'sd15;
	qsin_lut[5370] = -9'sd73;
	icos_lut[5370] =  9'sd30;
	qsin_lut[5371] = -9'sd66;
	icos_lut[5371] =  9'sd44;
	qsin_lut[5372] = -9'sd56;
	icos_lut[5372] =  9'sd56;
	qsin_lut[5373] = -9'sd44;
	icos_lut[5373] =  9'sd66;
	qsin_lut[5374] = -9'sd30;
	icos_lut[5374] =  9'sd73;
	qsin_lut[5375] = -9'sd15;
	icos_lut[5375] =  9'sd77;
	qsin_lut[5376] =  9'sd0;
	icos_lut[5376] =  9'sd81;
	qsin_lut[5377] =  9'sd16;
	icos_lut[5377] =  9'sd79;
	qsin_lut[5378] =  9'sd31;
	icos_lut[5378] =  9'sd75;
	qsin_lut[5379] =  9'sd45;
	icos_lut[5379] =  9'sd67;
	qsin_lut[5380] =  9'sd57;
	icos_lut[5380] =  9'sd57;
	qsin_lut[5381] =  9'sd67;
	icos_lut[5381] =  9'sd45;
	qsin_lut[5382] =  9'sd75;
	icos_lut[5382] =  9'sd31;
	qsin_lut[5383] =  9'sd79;
	icos_lut[5383] =  9'sd16;
	qsin_lut[5384] =  9'sd81;
	icos_lut[5384] =  9'sd0;
	qsin_lut[5385] =  9'sd79;
	icos_lut[5385] = -9'sd16;
	qsin_lut[5386] =  9'sd75;
	icos_lut[5386] = -9'sd31;
	qsin_lut[5387] =  9'sd67;
	icos_lut[5387] = -9'sd45;
	qsin_lut[5388] =  9'sd57;
	icos_lut[5388] = -9'sd57;
	qsin_lut[5389] =  9'sd45;
	icos_lut[5389] = -9'sd67;
	qsin_lut[5390] =  9'sd31;
	icos_lut[5390] = -9'sd75;
	qsin_lut[5391] =  9'sd16;
	icos_lut[5391] = -9'sd79;
	qsin_lut[5392] =  9'sd0;
	icos_lut[5392] = -9'sd81;
	qsin_lut[5393] = -9'sd16;
	icos_lut[5393] = -9'sd79;
	qsin_lut[5394] = -9'sd31;
	icos_lut[5394] = -9'sd75;
	qsin_lut[5395] = -9'sd45;
	icos_lut[5395] = -9'sd67;
	qsin_lut[5396] = -9'sd57;
	icos_lut[5396] = -9'sd57;
	qsin_lut[5397] = -9'sd67;
	icos_lut[5397] = -9'sd45;
	qsin_lut[5398] = -9'sd75;
	icos_lut[5398] = -9'sd31;
	qsin_lut[5399] = -9'sd79;
	icos_lut[5399] = -9'sd16;
	qsin_lut[5400] = -9'sd81;
	icos_lut[5400] = -9'sd0;
	qsin_lut[5401] = -9'sd79;
	icos_lut[5401] =  9'sd16;
	qsin_lut[5402] = -9'sd75;
	icos_lut[5402] =  9'sd31;
	qsin_lut[5403] = -9'sd67;
	icos_lut[5403] =  9'sd45;
	qsin_lut[5404] = -9'sd57;
	icos_lut[5404] =  9'sd57;
	qsin_lut[5405] = -9'sd45;
	icos_lut[5405] =  9'sd67;
	qsin_lut[5406] = -9'sd31;
	icos_lut[5406] =  9'sd75;
	qsin_lut[5407] = -9'sd16;
	icos_lut[5407] =  9'sd79;
	qsin_lut[5408] =  9'sd0;
	icos_lut[5408] =  9'sd83;
	qsin_lut[5409] =  9'sd16;
	icos_lut[5409] =  9'sd81;
	qsin_lut[5410] =  9'sd32;
	icos_lut[5410] =  9'sd77;
	qsin_lut[5411] =  9'sd46;
	icos_lut[5411] =  9'sd69;
	qsin_lut[5412] =  9'sd59;
	icos_lut[5412] =  9'sd59;
	qsin_lut[5413] =  9'sd69;
	icos_lut[5413] =  9'sd46;
	qsin_lut[5414] =  9'sd77;
	icos_lut[5414] =  9'sd32;
	qsin_lut[5415] =  9'sd81;
	icos_lut[5415] =  9'sd16;
	qsin_lut[5416] =  9'sd83;
	icos_lut[5416] =  9'sd0;
	qsin_lut[5417] =  9'sd81;
	icos_lut[5417] = -9'sd16;
	qsin_lut[5418] =  9'sd77;
	icos_lut[5418] = -9'sd32;
	qsin_lut[5419] =  9'sd69;
	icos_lut[5419] = -9'sd46;
	qsin_lut[5420] =  9'sd59;
	icos_lut[5420] = -9'sd59;
	qsin_lut[5421] =  9'sd46;
	icos_lut[5421] = -9'sd69;
	qsin_lut[5422] =  9'sd32;
	icos_lut[5422] = -9'sd77;
	qsin_lut[5423] =  9'sd16;
	icos_lut[5423] = -9'sd81;
	qsin_lut[5424] =  9'sd0;
	icos_lut[5424] = -9'sd83;
	qsin_lut[5425] = -9'sd16;
	icos_lut[5425] = -9'sd81;
	qsin_lut[5426] = -9'sd32;
	icos_lut[5426] = -9'sd77;
	qsin_lut[5427] = -9'sd46;
	icos_lut[5427] = -9'sd69;
	qsin_lut[5428] = -9'sd59;
	icos_lut[5428] = -9'sd59;
	qsin_lut[5429] = -9'sd69;
	icos_lut[5429] = -9'sd46;
	qsin_lut[5430] = -9'sd77;
	icos_lut[5430] = -9'sd32;
	qsin_lut[5431] = -9'sd81;
	icos_lut[5431] = -9'sd16;
	qsin_lut[5432] = -9'sd83;
	icos_lut[5432] = -9'sd0;
	qsin_lut[5433] = -9'sd81;
	icos_lut[5433] =  9'sd16;
	qsin_lut[5434] = -9'sd77;
	icos_lut[5434] =  9'sd32;
	qsin_lut[5435] = -9'sd69;
	icos_lut[5435] =  9'sd46;
	qsin_lut[5436] = -9'sd59;
	icos_lut[5436] =  9'sd59;
	qsin_lut[5437] = -9'sd46;
	icos_lut[5437] =  9'sd69;
	qsin_lut[5438] = -9'sd32;
	icos_lut[5438] =  9'sd77;
	qsin_lut[5439] = -9'sd16;
	icos_lut[5439] =  9'sd81;
	qsin_lut[5440] =  9'sd0;
	icos_lut[5440] =  9'sd85;
	qsin_lut[5441] =  9'sd17;
	icos_lut[5441] =  9'sd83;
	qsin_lut[5442] =  9'sd33;
	icos_lut[5442] =  9'sd79;
	qsin_lut[5443] =  9'sd47;
	icos_lut[5443] =  9'sd71;
	qsin_lut[5444] =  9'sd60;
	icos_lut[5444] =  9'sd60;
	qsin_lut[5445] =  9'sd71;
	icos_lut[5445] =  9'sd47;
	qsin_lut[5446] =  9'sd79;
	icos_lut[5446] =  9'sd33;
	qsin_lut[5447] =  9'sd83;
	icos_lut[5447] =  9'sd17;
	qsin_lut[5448] =  9'sd85;
	icos_lut[5448] =  9'sd0;
	qsin_lut[5449] =  9'sd83;
	icos_lut[5449] = -9'sd17;
	qsin_lut[5450] =  9'sd79;
	icos_lut[5450] = -9'sd33;
	qsin_lut[5451] =  9'sd71;
	icos_lut[5451] = -9'sd47;
	qsin_lut[5452] =  9'sd60;
	icos_lut[5452] = -9'sd60;
	qsin_lut[5453] =  9'sd47;
	icos_lut[5453] = -9'sd71;
	qsin_lut[5454] =  9'sd33;
	icos_lut[5454] = -9'sd79;
	qsin_lut[5455] =  9'sd17;
	icos_lut[5455] = -9'sd83;
	qsin_lut[5456] =  9'sd0;
	icos_lut[5456] = -9'sd85;
	qsin_lut[5457] = -9'sd17;
	icos_lut[5457] = -9'sd83;
	qsin_lut[5458] = -9'sd33;
	icos_lut[5458] = -9'sd79;
	qsin_lut[5459] = -9'sd47;
	icos_lut[5459] = -9'sd71;
	qsin_lut[5460] = -9'sd60;
	icos_lut[5460] = -9'sd60;
	qsin_lut[5461] = -9'sd71;
	icos_lut[5461] = -9'sd47;
	qsin_lut[5462] = -9'sd79;
	icos_lut[5462] = -9'sd33;
	qsin_lut[5463] = -9'sd83;
	icos_lut[5463] = -9'sd17;
	qsin_lut[5464] = -9'sd85;
	icos_lut[5464] = -9'sd0;
	qsin_lut[5465] = -9'sd83;
	icos_lut[5465] =  9'sd17;
	qsin_lut[5466] = -9'sd79;
	icos_lut[5466] =  9'sd33;
	qsin_lut[5467] = -9'sd71;
	icos_lut[5467] =  9'sd47;
	qsin_lut[5468] = -9'sd60;
	icos_lut[5468] =  9'sd60;
	qsin_lut[5469] = -9'sd47;
	icos_lut[5469] =  9'sd71;
	qsin_lut[5470] = -9'sd33;
	icos_lut[5470] =  9'sd79;
	qsin_lut[5471] = -9'sd17;
	icos_lut[5471] =  9'sd83;
	qsin_lut[5472] =  9'sd0;
	icos_lut[5472] =  9'sd87;
	qsin_lut[5473] =  9'sd17;
	icos_lut[5473] =  9'sd85;
	qsin_lut[5474] =  9'sd33;
	icos_lut[5474] =  9'sd80;
	qsin_lut[5475] =  9'sd48;
	icos_lut[5475] =  9'sd72;
	qsin_lut[5476] =  9'sd62;
	icos_lut[5476] =  9'sd62;
	qsin_lut[5477] =  9'sd72;
	icos_lut[5477] =  9'sd48;
	qsin_lut[5478] =  9'sd80;
	icos_lut[5478] =  9'sd33;
	qsin_lut[5479] =  9'sd85;
	icos_lut[5479] =  9'sd17;
	qsin_lut[5480] =  9'sd87;
	icos_lut[5480] =  9'sd0;
	qsin_lut[5481] =  9'sd85;
	icos_lut[5481] = -9'sd17;
	qsin_lut[5482] =  9'sd80;
	icos_lut[5482] = -9'sd33;
	qsin_lut[5483] =  9'sd72;
	icos_lut[5483] = -9'sd48;
	qsin_lut[5484] =  9'sd62;
	icos_lut[5484] = -9'sd62;
	qsin_lut[5485] =  9'sd48;
	icos_lut[5485] = -9'sd72;
	qsin_lut[5486] =  9'sd33;
	icos_lut[5486] = -9'sd80;
	qsin_lut[5487] =  9'sd17;
	icos_lut[5487] = -9'sd85;
	qsin_lut[5488] =  9'sd0;
	icos_lut[5488] = -9'sd87;
	qsin_lut[5489] = -9'sd17;
	icos_lut[5489] = -9'sd85;
	qsin_lut[5490] = -9'sd33;
	icos_lut[5490] = -9'sd80;
	qsin_lut[5491] = -9'sd48;
	icos_lut[5491] = -9'sd72;
	qsin_lut[5492] = -9'sd62;
	icos_lut[5492] = -9'sd62;
	qsin_lut[5493] = -9'sd72;
	icos_lut[5493] = -9'sd48;
	qsin_lut[5494] = -9'sd80;
	icos_lut[5494] = -9'sd33;
	qsin_lut[5495] = -9'sd85;
	icos_lut[5495] = -9'sd17;
	qsin_lut[5496] = -9'sd87;
	icos_lut[5496] = -9'sd0;
	qsin_lut[5497] = -9'sd85;
	icos_lut[5497] =  9'sd17;
	qsin_lut[5498] = -9'sd80;
	icos_lut[5498] =  9'sd33;
	qsin_lut[5499] = -9'sd72;
	icos_lut[5499] =  9'sd48;
	qsin_lut[5500] = -9'sd62;
	icos_lut[5500] =  9'sd62;
	qsin_lut[5501] = -9'sd48;
	icos_lut[5501] =  9'sd72;
	qsin_lut[5502] = -9'sd33;
	icos_lut[5502] =  9'sd80;
	qsin_lut[5503] = -9'sd17;
	icos_lut[5503] =  9'sd85;
	qsin_lut[5504] =  9'sd0;
	icos_lut[5504] =  9'sd89;
	qsin_lut[5505] =  9'sd17;
	icos_lut[5505] =  9'sd87;
	qsin_lut[5506] =  9'sd34;
	icos_lut[5506] =  9'sd82;
	qsin_lut[5507] =  9'sd49;
	icos_lut[5507] =  9'sd74;
	qsin_lut[5508] =  9'sd63;
	icos_lut[5508] =  9'sd63;
	qsin_lut[5509] =  9'sd74;
	icos_lut[5509] =  9'sd49;
	qsin_lut[5510] =  9'sd82;
	icos_lut[5510] =  9'sd34;
	qsin_lut[5511] =  9'sd87;
	icos_lut[5511] =  9'sd17;
	qsin_lut[5512] =  9'sd89;
	icos_lut[5512] =  9'sd0;
	qsin_lut[5513] =  9'sd87;
	icos_lut[5513] = -9'sd17;
	qsin_lut[5514] =  9'sd82;
	icos_lut[5514] = -9'sd34;
	qsin_lut[5515] =  9'sd74;
	icos_lut[5515] = -9'sd49;
	qsin_lut[5516] =  9'sd63;
	icos_lut[5516] = -9'sd63;
	qsin_lut[5517] =  9'sd49;
	icos_lut[5517] = -9'sd74;
	qsin_lut[5518] =  9'sd34;
	icos_lut[5518] = -9'sd82;
	qsin_lut[5519] =  9'sd17;
	icos_lut[5519] = -9'sd87;
	qsin_lut[5520] =  9'sd0;
	icos_lut[5520] = -9'sd89;
	qsin_lut[5521] = -9'sd17;
	icos_lut[5521] = -9'sd87;
	qsin_lut[5522] = -9'sd34;
	icos_lut[5522] = -9'sd82;
	qsin_lut[5523] = -9'sd49;
	icos_lut[5523] = -9'sd74;
	qsin_lut[5524] = -9'sd63;
	icos_lut[5524] = -9'sd63;
	qsin_lut[5525] = -9'sd74;
	icos_lut[5525] = -9'sd49;
	qsin_lut[5526] = -9'sd82;
	icos_lut[5526] = -9'sd34;
	qsin_lut[5527] = -9'sd87;
	icos_lut[5527] = -9'sd17;
	qsin_lut[5528] = -9'sd89;
	icos_lut[5528] = -9'sd0;
	qsin_lut[5529] = -9'sd87;
	icos_lut[5529] =  9'sd17;
	qsin_lut[5530] = -9'sd82;
	icos_lut[5530] =  9'sd34;
	qsin_lut[5531] = -9'sd74;
	icos_lut[5531] =  9'sd49;
	qsin_lut[5532] = -9'sd63;
	icos_lut[5532] =  9'sd63;
	qsin_lut[5533] = -9'sd49;
	icos_lut[5533] =  9'sd74;
	qsin_lut[5534] = -9'sd34;
	icos_lut[5534] =  9'sd82;
	qsin_lut[5535] = -9'sd17;
	icos_lut[5535] =  9'sd87;
	qsin_lut[5536] =  9'sd0;
	icos_lut[5536] =  9'sd91;
	qsin_lut[5537] =  9'sd18;
	icos_lut[5537] =  9'sd89;
	qsin_lut[5538] =  9'sd35;
	icos_lut[5538] =  9'sd84;
	qsin_lut[5539] =  9'sd51;
	icos_lut[5539] =  9'sd76;
	qsin_lut[5540] =  9'sd64;
	icos_lut[5540] =  9'sd64;
	qsin_lut[5541] =  9'sd76;
	icos_lut[5541] =  9'sd51;
	qsin_lut[5542] =  9'sd84;
	icos_lut[5542] =  9'sd35;
	qsin_lut[5543] =  9'sd89;
	icos_lut[5543] =  9'sd18;
	qsin_lut[5544] =  9'sd91;
	icos_lut[5544] =  9'sd0;
	qsin_lut[5545] =  9'sd89;
	icos_lut[5545] = -9'sd18;
	qsin_lut[5546] =  9'sd84;
	icos_lut[5546] = -9'sd35;
	qsin_lut[5547] =  9'sd76;
	icos_lut[5547] = -9'sd51;
	qsin_lut[5548] =  9'sd64;
	icos_lut[5548] = -9'sd64;
	qsin_lut[5549] =  9'sd51;
	icos_lut[5549] = -9'sd76;
	qsin_lut[5550] =  9'sd35;
	icos_lut[5550] = -9'sd84;
	qsin_lut[5551] =  9'sd18;
	icos_lut[5551] = -9'sd89;
	qsin_lut[5552] =  9'sd0;
	icos_lut[5552] = -9'sd91;
	qsin_lut[5553] = -9'sd18;
	icos_lut[5553] = -9'sd89;
	qsin_lut[5554] = -9'sd35;
	icos_lut[5554] = -9'sd84;
	qsin_lut[5555] = -9'sd51;
	icos_lut[5555] = -9'sd76;
	qsin_lut[5556] = -9'sd64;
	icos_lut[5556] = -9'sd64;
	qsin_lut[5557] = -9'sd76;
	icos_lut[5557] = -9'sd51;
	qsin_lut[5558] = -9'sd84;
	icos_lut[5558] = -9'sd35;
	qsin_lut[5559] = -9'sd89;
	icos_lut[5559] = -9'sd18;
	qsin_lut[5560] = -9'sd91;
	icos_lut[5560] = -9'sd0;
	qsin_lut[5561] = -9'sd89;
	icos_lut[5561] =  9'sd18;
	qsin_lut[5562] = -9'sd84;
	icos_lut[5562] =  9'sd35;
	qsin_lut[5563] = -9'sd76;
	icos_lut[5563] =  9'sd51;
	qsin_lut[5564] = -9'sd64;
	icos_lut[5564] =  9'sd64;
	qsin_lut[5565] = -9'sd51;
	icos_lut[5565] =  9'sd76;
	qsin_lut[5566] = -9'sd35;
	icos_lut[5566] =  9'sd84;
	qsin_lut[5567] = -9'sd18;
	icos_lut[5567] =  9'sd89;
	qsin_lut[5568] =  9'sd0;
	icos_lut[5568] =  9'sd93;
	qsin_lut[5569] =  9'sd18;
	icos_lut[5569] =  9'sd91;
	qsin_lut[5570] =  9'sd36;
	icos_lut[5570] =  9'sd86;
	qsin_lut[5571] =  9'sd52;
	icos_lut[5571] =  9'sd77;
	qsin_lut[5572] =  9'sd66;
	icos_lut[5572] =  9'sd66;
	qsin_lut[5573] =  9'sd77;
	icos_lut[5573] =  9'sd52;
	qsin_lut[5574] =  9'sd86;
	icos_lut[5574] =  9'sd36;
	qsin_lut[5575] =  9'sd91;
	icos_lut[5575] =  9'sd18;
	qsin_lut[5576] =  9'sd93;
	icos_lut[5576] =  9'sd0;
	qsin_lut[5577] =  9'sd91;
	icos_lut[5577] = -9'sd18;
	qsin_lut[5578] =  9'sd86;
	icos_lut[5578] = -9'sd36;
	qsin_lut[5579] =  9'sd77;
	icos_lut[5579] = -9'sd52;
	qsin_lut[5580] =  9'sd66;
	icos_lut[5580] = -9'sd66;
	qsin_lut[5581] =  9'sd52;
	icos_lut[5581] = -9'sd77;
	qsin_lut[5582] =  9'sd36;
	icos_lut[5582] = -9'sd86;
	qsin_lut[5583] =  9'sd18;
	icos_lut[5583] = -9'sd91;
	qsin_lut[5584] =  9'sd0;
	icos_lut[5584] = -9'sd93;
	qsin_lut[5585] = -9'sd18;
	icos_lut[5585] = -9'sd91;
	qsin_lut[5586] = -9'sd36;
	icos_lut[5586] = -9'sd86;
	qsin_lut[5587] = -9'sd52;
	icos_lut[5587] = -9'sd77;
	qsin_lut[5588] = -9'sd66;
	icos_lut[5588] = -9'sd66;
	qsin_lut[5589] = -9'sd77;
	icos_lut[5589] = -9'sd52;
	qsin_lut[5590] = -9'sd86;
	icos_lut[5590] = -9'sd36;
	qsin_lut[5591] = -9'sd91;
	icos_lut[5591] = -9'sd18;
	qsin_lut[5592] = -9'sd93;
	icos_lut[5592] = -9'sd0;
	qsin_lut[5593] = -9'sd91;
	icos_lut[5593] =  9'sd18;
	qsin_lut[5594] = -9'sd86;
	icos_lut[5594] =  9'sd36;
	qsin_lut[5595] = -9'sd77;
	icos_lut[5595] =  9'sd52;
	qsin_lut[5596] = -9'sd66;
	icos_lut[5596] =  9'sd66;
	qsin_lut[5597] = -9'sd52;
	icos_lut[5597] =  9'sd77;
	qsin_lut[5598] = -9'sd36;
	icos_lut[5598] =  9'sd86;
	qsin_lut[5599] = -9'sd18;
	icos_lut[5599] =  9'sd91;
	qsin_lut[5600] =  9'sd0;
	icos_lut[5600] =  9'sd95;
	qsin_lut[5601] =  9'sd19;
	icos_lut[5601] =  9'sd93;
	qsin_lut[5602] =  9'sd36;
	icos_lut[5602] =  9'sd88;
	qsin_lut[5603] =  9'sd53;
	icos_lut[5603] =  9'sd79;
	qsin_lut[5604] =  9'sd67;
	icos_lut[5604] =  9'sd67;
	qsin_lut[5605] =  9'sd79;
	icos_lut[5605] =  9'sd53;
	qsin_lut[5606] =  9'sd88;
	icos_lut[5606] =  9'sd36;
	qsin_lut[5607] =  9'sd93;
	icos_lut[5607] =  9'sd19;
	qsin_lut[5608] =  9'sd95;
	icos_lut[5608] =  9'sd0;
	qsin_lut[5609] =  9'sd93;
	icos_lut[5609] = -9'sd19;
	qsin_lut[5610] =  9'sd88;
	icos_lut[5610] = -9'sd36;
	qsin_lut[5611] =  9'sd79;
	icos_lut[5611] = -9'sd53;
	qsin_lut[5612] =  9'sd67;
	icos_lut[5612] = -9'sd67;
	qsin_lut[5613] =  9'sd53;
	icos_lut[5613] = -9'sd79;
	qsin_lut[5614] =  9'sd36;
	icos_lut[5614] = -9'sd88;
	qsin_lut[5615] =  9'sd19;
	icos_lut[5615] = -9'sd93;
	qsin_lut[5616] =  9'sd0;
	icos_lut[5616] = -9'sd95;
	qsin_lut[5617] = -9'sd19;
	icos_lut[5617] = -9'sd93;
	qsin_lut[5618] = -9'sd36;
	icos_lut[5618] = -9'sd88;
	qsin_lut[5619] = -9'sd53;
	icos_lut[5619] = -9'sd79;
	qsin_lut[5620] = -9'sd67;
	icos_lut[5620] = -9'sd67;
	qsin_lut[5621] = -9'sd79;
	icos_lut[5621] = -9'sd53;
	qsin_lut[5622] = -9'sd88;
	icos_lut[5622] = -9'sd36;
	qsin_lut[5623] = -9'sd93;
	icos_lut[5623] = -9'sd19;
	qsin_lut[5624] = -9'sd95;
	icos_lut[5624] = -9'sd0;
	qsin_lut[5625] = -9'sd93;
	icos_lut[5625] =  9'sd19;
	qsin_lut[5626] = -9'sd88;
	icos_lut[5626] =  9'sd36;
	qsin_lut[5627] = -9'sd79;
	icos_lut[5627] =  9'sd53;
	qsin_lut[5628] = -9'sd67;
	icos_lut[5628] =  9'sd67;
	qsin_lut[5629] = -9'sd53;
	icos_lut[5629] =  9'sd79;
	qsin_lut[5630] = -9'sd36;
	icos_lut[5630] =  9'sd88;
	qsin_lut[5631] = -9'sd19;
	icos_lut[5631] =  9'sd93;
	qsin_lut[5632] =  9'sd0;
	icos_lut[5632] =  9'sd97;
	qsin_lut[5633] =  9'sd19;
	icos_lut[5633] =  9'sd95;
	qsin_lut[5634] =  9'sd37;
	icos_lut[5634] =  9'sd90;
	qsin_lut[5635] =  9'sd54;
	icos_lut[5635] =  9'sd81;
	qsin_lut[5636] =  9'sd69;
	icos_lut[5636] =  9'sd69;
	qsin_lut[5637] =  9'sd81;
	icos_lut[5637] =  9'sd54;
	qsin_lut[5638] =  9'sd90;
	icos_lut[5638] =  9'sd37;
	qsin_lut[5639] =  9'sd95;
	icos_lut[5639] =  9'sd19;
	qsin_lut[5640] =  9'sd97;
	icos_lut[5640] =  9'sd0;
	qsin_lut[5641] =  9'sd95;
	icos_lut[5641] = -9'sd19;
	qsin_lut[5642] =  9'sd90;
	icos_lut[5642] = -9'sd37;
	qsin_lut[5643] =  9'sd81;
	icos_lut[5643] = -9'sd54;
	qsin_lut[5644] =  9'sd69;
	icos_lut[5644] = -9'sd69;
	qsin_lut[5645] =  9'sd54;
	icos_lut[5645] = -9'sd81;
	qsin_lut[5646] =  9'sd37;
	icos_lut[5646] = -9'sd90;
	qsin_lut[5647] =  9'sd19;
	icos_lut[5647] = -9'sd95;
	qsin_lut[5648] =  9'sd0;
	icos_lut[5648] = -9'sd97;
	qsin_lut[5649] = -9'sd19;
	icos_lut[5649] = -9'sd95;
	qsin_lut[5650] = -9'sd37;
	icos_lut[5650] = -9'sd90;
	qsin_lut[5651] = -9'sd54;
	icos_lut[5651] = -9'sd81;
	qsin_lut[5652] = -9'sd69;
	icos_lut[5652] = -9'sd69;
	qsin_lut[5653] = -9'sd81;
	icos_lut[5653] = -9'sd54;
	qsin_lut[5654] = -9'sd90;
	icos_lut[5654] = -9'sd37;
	qsin_lut[5655] = -9'sd95;
	icos_lut[5655] = -9'sd19;
	qsin_lut[5656] = -9'sd97;
	icos_lut[5656] = -9'sd0;
	qsin_lut[5657] = -9'sd95;
	icos_lut[5657] =  9'sd19;
	qsin_lut[5658] = -9'sd90;
	icos_lut[5658] =  9'sd37;
	qsin_lut[5659] = -9'sd81;
	icos_lut[5659] =  9'sd54;
	qsin_lut[5660] = -9'sd69;
	icos_lut[5660] =  9'sd69;
	qsin_lut[5661] = -9'sd54;
	icos_lut[5661] =  9'sd81;
	qsin_lut[5662] = -9'sd37;
	icos_lut[5662] =  9'sd90;
	qsin_lut[5663] = -9'sd19;
	icos_lut[5663] =  9'sd95;
	qsin_lut[5664] =  9'sd0;
	icos_lut[5664] =  9'sd99;
	qsin_lut[5665] =  9'sd19;
	icos_lut[5665] =  9'sd97;
	qsin_lut[5666] =  9'sd38;
	icos_lut[5666] =  9'sd91;
	qsin_lut[5667] =  9'sd55;
	icos_lut[5667] =  9'sd82;
	qsin_lut[5668] =  9'sd70;
	icos_lut[5668] =  9'sd70;
	qsin_lut[5669] =  9'sd82;
	icos_lut[5669] =  9'sd55;
	qsin_lut[5670] =  9'sd91;
	icos_lut[5670] =  9'sd38;
	qsin_lut[5671] =  9'sd97;
	icos_lut[5671] =  9'sd19;
	qsin_lut[5672] =  9'sd99;
	icos_lut[5672] =  9'sd0;
	qsin_lut[5673] =  9'sd97;
	icos_lut[5673] = -9'sd19;
	qsin_lut[5674] =  9'sd91;
	icos_lut[5674] = -9'sd38;
	qsin_lut[5675] =  9'sd82;
	icos_lut[5675] = -9'sd55;
	qsin_lut[5676] =  9'sd70;
	icos_lut[5676] = -9'sd70;
	qsin_lut[5677] =  9'sd55;
	icos_lut[5677] = -9'sd82;
	qsin_lut[5678] =  9'sd38;
	icos_lut[5678] = -9'sd91;
	qsin_lut[5679] =  9'sd19;
	icos_lut[5679] = -9'sd97;
	qsin_lut[5680] =  9'sd0;
	icos_lut[5680] = -9'sd99;
	qsin_lut[5681] = -9'sd19;
	icos_lut[5681] = -9'sd97;
	qsin_lut[5682] = -9'sd38;
	icos_lut[5682] = -9'sd91;
	qsin_lut[5683] = -9'sd55;
	icos_lut[5683] = -9'sd82;
	qsin_lut[5684] = -9'sd70;
	icos_lut[5684] = -9'sd70;
	qsin_lut[5685] = -9'sd82;
	icos_lut[5685] = -9'sd55;
	qsin_lut[5686] = -9'sd91;
	icos_lut[5686] = -9'sd38;
	qsin_lut[5687] = -9'sd97;
	icos_lut[5687] = -9'sd19;
	qsin_lut[5688] = -9'sd99;
	icos_lut[5688] = -9'sd0;
	qsin_lut[5689] = -9'sd97;
	icos_lut[5689] =  9'sd19;
	qsin_lut[5690] = -9'sd91;
	icos_lut[5690] =  9'sd38;
	qsin_lut[5691] = -9'sd82;
	icos_lut[5691] =  9'sd55;
	qsin_lut[5692] = -9'sd70;
	icos_lut[5692] =  9'sd70;
	qsin_lut[5693] = -9'sd55;
	icos_lut[5693] =  9'sd82;
	qsin_lut[5694] = -9'sd38;
	icos_lut[5694] =  9'sd91;
	qsin_lut[5695] = -9'sd19;
	icos_lut[5695] =  9'sd97;
	qsin_lut[5696] =  9'sd0;
	icos_lut[5696] =  9'sd101;
	qsin_lut[5697] =  9'sd20;
	icos_lut[5697] =  9'sd99;
	qsin_lut[5698] =  9'sd39;
	icos_lut[5698] =  9'sd93;
	qsin_lut[5699] =  9'sd56;
	icos_lut[5699] =  9'sd84;
	qsin_lut[5700] =  9'sd71;
	icos_lut[5700] =  9'sd71;
	qsin_lut[5701] =  9'sd84;
	icos_lut[5701] =  9'sd56;
	qsin_lut[5702] =  9'sd93;
	icos_lut[5702] =  9'sd39;
	qsin_lut[5703] =  9'sd99;
	icos_lut[5703] =  9'sd20;
	qsin_lut[5704] =  9'sd101;
	icos_lut[5704] =  9'sd0;
	qsin_lut[5705] =  9'sd99;
	icos_lut[5705] = -9'sd20;
	qsin_lut[5706] =  9'sd93;
	icos_lut[5706] = -9'sd39;
	qsin_lut[5707] =  9'sd84;
	icos_lut[5707] = -9'sd56;
	qsin_lut[5708] =  9'sd71;
	icos_lut[5708] = -9'sd71;
	qsin_lut[5709] =  9'sd56;
	icos_lut[5709] = -9'sd84;
	qsin_lut[5710] =  9'sd39;
	icos_lut[5710] = -9'sd93;
	qsin_lut[5711] =  9'sd20;
	icos_lut[5711] = -9'sd99;
	qsin_lut[5712] =  9'sd0;
	icos_lut[5712] = -9'sd101;
	qsin_lut[5713] = -9'sd20;
	icos_lut[5713] = -9'sd99;
	qsin_lut[5714] = -9'sd39;
	icos_lut[5714] = -9'sd93;
	qsin_lut[5715] = -9'sd56;
	icos_lut[5715] = -9'sd84;
	qsin_lut[5716] = -9'sd71;
	icos_lut[5716] = -9'sd71;
	qsin_lut[5717] = -9'sd84;
	icos_lut[5717] = -9'sd56;
	qsin_lut[5718] = -9'sd93;
	icos_lut[5718] = -9'sd39;
	qsin_lut[5719] = -9'sd99;
	icos_lut[5719] = -9'sd20;
	qsin_lut[5720] = -9'sd101;
	icos_lut[5720] = -9'sd0;
	qsin_lut[5721] = -9'sd99;
	icos_lut[5721] =  9'sd20;
	qsin_lut[5722] = -9'sd93;
	icos_lut[5722] =  9'sd39;
	qsin_lut[5723] = -9'sd84;
	icos_lut[5723] =  9'sd56;
	qsin_lut[5724] = -9'sd71;
	icos_lut[5724] =  9'sd71;
	qsin_lut[5725] = -9'sd56;
	icos_lut[5725] =  9'sd84;
	qsin_lut[5726] = -9'sd39;
	icos_lut[5726] =  9'sd93;
	qsin_lut[5727] = -9'sd20;
	icos_lut[5727] =  9'sd99;
	qsin_lut[5728] =  9'sd0;
	icos_lut[5728] =  9'sd103;
	qsin_lut[5729] =  9'sd20;
	icos_lut[5729] =  9'sd101;
	qsin_lut[5730] =  9'sd39;
	icos_lut[5730] =  9'sd95;
	qsin_lut[5731] =  9'sd57;
	icos_lut[5731] =  9'sd86;
	qsin_lut[5732] =  9'sd73;
	icos_lut[5732] =  9'sd73;
	qsin_lut[5733] =  9'sd86;
	icos_lut[5733] =  9'sd57;
	qsin_lut[5734] =  9'sd95;
	icos_lut[5734] =  9'sd39;
	qsin_lut[5735] =  9'sd101;
	icos_lut[5735] =  9'sd20;
	qsin_lut[5736] =  9'sd103;
	icos_lut[5736] =  9'sd0;
	qsin_lut[5737] =  9'sd101;
	icos_lut[5737] = -9'sd20;
	qsin_lut[5738] =  9'sd95;
	icos_lut[5738] = -9'sd39;
	qsin_lut[5739] =  9'sd86;
	icos_lut[5739] = -9'sd57;
	qsin_lut[5740] =  9'sd73;
	icos_lut[5740] = -9'sd73;
	qsin_lut[5741] =  9'sd57;
	icos_lut[5741] = -9'sd86;
	qsin_lut[5742] =  9'sd39;
	icos_lut[5742] = -9'sd95;
	qsin_lut[5743] =  9'sd20;
	icos_lut[5743] = -9'sd101;
	qsin_lut[5744] =  9'sd0;
	icos_lut[5744] = -9'sd103;
	qsin_lut[5745] = -9'sd20;
	icos_lut[5745] = -9'sd101;
	qsin_lut[5746] = -9'sd39;
	icos_lut[5746] = -9'sd95;
	qsin_lut[5747] = -9'sd57;
	icos_lut[5747] = -9'sd86;
	qsin_lut[5748] = -9'sd73;
	icos_lut[5748] = -9'sd73;
	qsin_lut[5749] = -9'sd86;
	icos_lut[5749] = -9'sd57;
	qsin_lut[5750] = -9'sd95;
	icos_lut[5750] = -9'sd39;
	qsin_lut[5751] = -9'sd101;
	icos_lut[5751] = -9'sd20;
	qsin_lut[5752] = -9'sd103;
	icos_lut[5752] = -9'sd0;
	qsin_lut[5753] = -9'sd101;
	icos_lut[5753] =  9'sd20;
	qsin_lut[5754] = -9'sd95;
	icos_lut[5754] =  9'sd39;
	qsin_lut[5755] = -9'sd86;
	icos_lut[5755] =  9'sd57;
	qsin_lut[5756] = -9'sd73;
	icos_lut[5756] =  9'sd73;
	qsin_lut[5757] = -9'sd57;
	icos_lut[5757] =  9'sd86;
	qsin_lut[5758] = -9'sd39;
	icos_lut[5758] =  9'sd95;
	qsin_lut[5759] = -9'sd20;
	icos_lut[5759] =  9'sd101;
	qsin_lut[5760] =  9'sd0;
	icos_lut[5760] =  9'sd105;
	qsin_lut[5761] =  9'sd20;
	icos_lut[5761] =  9'sd103;
	qsin_lut[5762] =  9'sd40;
	icos_lut[5762] =  9'sd97;
	qsin_lut[5763] =  9'sd58;
	icos_lut[5763] =  9'sd87;
	qsin_lut[5764] =  9'sd74;
	icos_lut[5764] =  9'sd74;
	qsin_lut[5765] =  9'sd87;
	icos_lut[5765] =  9'sd58;
	qsin_lut[5766] =  9'sd97;
	icos_lut[5766] =  9'sd40;
	qsin_lut[5767] =  9'sd103;
	icos_lut[5767] =  9'sd20;
	qsin_lut[5768] =  9'sd105;
	icos_lut[5768] =  9'sd0;
	qsin_lut[5769] =  9'sd103;
	icos_lut[5769] = -9'sd20;
	qsin_lut[5770] =  9'sd97;
	icos_lut[5770] = -9'sd40;
	qsin_lut[5771] =  9'sd87;
	icos_lut[5771] = -9'sd58;
	qsin_lut[5772] =  9'sd74;
	icos_lut[5772] = -9'sd74;
	qsin_lut[5773] =  9'sd58;
	icos_lut[5773] = -9'sd87;
	qsin_lut[5774] =  9'sd40;
	icos_lut[5774] = -9'sd97;
	qsin_lut[5775] =  9'sd20;
	icos_lut[5775] = -9'sd103;
	qsin_lut[5776] =  9'sd0;
	icos_lut[5776] = -9'sd105;
	qsin_lut[5777] = -9'sd20;
	icos_lut[5777] = -9'sd103;
	qsin_lut[5778] = -9'sd40;
	icos_lut[5778] = -9'sd97;
	qsin_lut[5779] = -9'sd58;
	icos_lut[5779] = -9'sd87;
	qsin_lut[5780] = -9'sd74;
	icos_lut[5780] = -9'sd74;
	qsin_lut[5781] = -9'sd87;
	icos_lut[5781] = -9'sd58;
	qsin_lut[5782] = -9'sd97;
	icos_lut[5782] = -9'sd40;
	qsin_lut[5783] = -9'sd103;
	icos_lut[5783] = -9'sd20;
	qsin_lut[5784] = -9'sd105;
	icos_lut[5784] = -9'sd0;
	qsin_lut[5785] = -9'sd103;
	icos_lut[5785] =  9'sd20;
	qsin_lut[5786] = -9'sd97;
	icos_lut[5786] =  9'sd40;
	qsin_lut[5787] = -9'sd87;
	icos_lut[5787] =  9'sd58;
	qsin_lut[5788] = -9'sd74;
	icos_lut[5788] =  9'sd74;
	qsin_lut[5789] = -9'sd58;
	icos_lut[5789] =  9'sd87;
	qsin_lut[5790] = -9'sd40;
	icos_lut[5790] =  9'sd97;
	qsin_lut[5791] = -9'sd20;
	icos_lut[5791] =  9'sd103;
	qsin_lut[5792] =  9'sd0;
	icos_lut[5792] =  9'sd107;
	qsin_lut[5793] =  9'sd21;
	icos_lut[5793] =  9'sd105;
	qsin_lut[5794] =  9'sd41;
	icos_lut[5794] =  9'sd99;
	qsin_lut[5795] =  9'sd59;
	icos_lut[5795] =  9'sd89;
	qsin_lut[5796] =  9'sd76;
	icos_lut[5796] =  9'sd76;
	qsin_lut[5797] =  9'sd89;
	icos_lut[5797] =  9'sd59;
	qsin_lut[5798] =  9'sd99;
	icos_lut[5798] =  9'sd41;
	qsin_lut[5799] =  9'sd105;
	icos_lut[5799] =  9'sd21;
	qsin_lut[5800] =  9'sd107;
	icos_lut[5800] =  9'sd0;
	qsin_lut[5801] =  9'sd105;
	icos_lut[5801] = -9'sd21;
	qsin_lut[5802] =  9'sd99;
	icos_lut[5802] = -9'sd41;
	qsin_lut[5803] =  9'sd89;
	icos_lut[5803] = -9'sd59;
	qsin_lut[5804] =  9'sd76;
	icos_lut[5804] = -9'sd76;
	qsin_lut[5805] =  9'sd59;
	icos_lut[5805] = -9'sd89;
	qsin_lut[5806] =  9'sd41;
	icos_lut[5806] = -9'sd99;
	qsin_lut[5807] =  9'sd21;
	icos_lut[5807] = -9'sd105;
	qsin_lut[5808] =  9'sd0;
	icos_lut[5808] = -9'sd107;
	qsin_lut[5809] = -9'sd21;
	icos_lut[5809] = -9'sd105;
	qsin_lut[5810] = -9'sd41;
	icos_lut[5810] = -9'sd99;
	qsin_lut[5811] = -9'sd59;
	icos_lut[5811] = -9'sd89;
	qsin_lut[5812] = -9'sd76;
	icos_lut[5812] = -9'sd76;
	qsin_lut[5813] = -9'sd89;
	icos_lut[5813] = -9'sd59;
	qsin_lut[5814] = -9'sd99;
	icos_lut[5814] = -9'sd41;
	qsin_lut[5815] = -9'sd105;
	icos_lut[5815] = -9'sd21;
	qsin_lut[5816] = -9'sd107;
	icos_lut[5816] = -9'sd0;
	qsin_lut[5817] = -9'sd105;
	icos_lut[5817] =  9'sd21;
	qsin_lut[5818] = -9'sd99;
	icos_lut[5818] =  9'sd41;
	qsin_lut[5819] = -9'sd89;
	icos_lut[5819] =  9'sd59;
	qsin_lut[5820] = -9'sd76;
	icos_lut[5820] =  9'sd76;
	qsin_lut[5821] = -9'sd59;
	icos_lut[5821] =  9'sd89;
	qsin_lut[5822] = -9'sd41;
	icos_lut[5822] =  9'sd99;
	qsin_lut[5823] = -9'sd21;
	icos_lut[5823] =  9'sd105;
	qsin_lut[5824] =  9'sd0;
	icos_lut[5824] =  9'sd109;
	qsin_lut[5825] =  9'sd21;
	icos_lut[5825] =  9'sd107;
	qsin_lut[5826] =  9'sd42;
	icos_lut[5826] =  9'sd101;
	qsin_lut[5827] =  9'sd61;
	icos_lut[5827] =  9'sd91;
	qsin_lut[5828] =  9'sd77;
	icos_lut[5828] =  9'sd77;
	qsin_lut[5829] =  9'sd91;
	icos_lut[5829] =  9'sd61;
	qsin_lut[5830] =  9'sd101;
	icos_lut[5830] =  9'sd42;
	qsin_lut[5831] =  9'sd107;
	icos_lut[5831] =  9'sd21;
	qsin_lut[5832] =  9'sd109;
	icos_lut[5832] =  9'sd0;
	qsin_lut[5833] =  9'sd107;
	icos_lut[5833] = -9'sd21;
	qsin_lut[5834] =  9'sd101;
	icos_lut[5834] = -9'sd42;
	qsin_lut[5835] =  9'sd91;
	icos_lut[5835] = -9'sd61;
	qsin_lut[5836] =  9'sd77;
	icos_lut[5836] = -9'sd77;
	qsin_lut[5837] =  9'sd61;
	icos_lut[5837] = -9'sd91;
	qsin_lut[5838] =  9'sd42;
	icos_lut[5838] = -9'sd101;
	qsin_lut[5839] =  9'sd21;
	icos_lut[5839] = -9'sd107;
	qsin_lut[5840] =  9'sd0;
	icos_lut[5840] = -9'sd109;
	qsin_lut[5841] = -9'sd21;
	icos_lut[5841] = -9'sd107;
	qsin_lut[5842] = -9'sd42;
	icos_lut[5842] = -9'sd101;
	qsin_lut[5843] = -9'sd61;
	icos_lut[5843] = -9'sd91;
	qsin_lut[5844] = -9'sd77;
	icos_lut[5844] = -9'sd77;
	qsin_lut[5845] = -9'sd91;
	icos_lut[5845] = -9'sd61;
	qsin_lut[5846] = -9'sd101;
	icos_lut[5846] = -9'sd42;
	qsin_lut[5847] = -9'sd107;
	icos_lut[5847] = -9'sd21;
	qsin_lut[5848] = -9'sd109;
	icos_lut[5848] = -9'sd0;
	qsin_lut[5849] = -9'sd107;
	icos_lut[5849] =  9'sd21;
	qsin_lut[5850] = -9'sd101;
	icos_lut[5850] =  9'sd42;
	qsin_lut[5851] = -9'sd91;
	icos_lut[5851] =  9'sd61;
	qsin_lut[5852] = -9'sd77;
	icos_lut[5852] =  9'sd77;
	qsin_lut[5853] = -9'sd61;
	icos_lut[5853] =  9'sd91;
	qsin_lut[5854] = -9'sd42;
	icos_lut[5854] =  9'sd101;
	qsin_lut[5855] = -9'sd21;
	icos_lut[5855] =  9'sd107;
	qsin_lut[5856] =  9'sd0;
	icos_lut[5856] =  9'sd111;
	qsin_lut[5857] =  9'sd22;
	icos_lut[5857] =  9'sd109;
	qsin_lut[5858] =  9'sd42;
	icos_lut[5858] =  9'sd103;
	qsin_lut[5859] =  9'sd62;
	icos_lut[5859] =  9'sd92;
	qsin_lut[5860] =  9'sd78;
	icos_lut[5860] =  9'sd78;
	qsin_lut[5861] =  9'sd92;
	icos_lut[5861] =  9'sd62;
	qsin_lut[5862] =  9'sd103;
	icos_lut[5862] =  9'sd42;
	qsin_lut[5863] =  9'sd109;
	icos_lut[5863] =  9'sd22;
	qsin_lut[5864] =  9'sd111;
	icos_lut[5864] =  9'sd0;
	qsin_lut[5865] =  9'sd109;
	icos_lut[5865] = -9'sd22;
	qsin_lut[5866] =  9'sd103;
	icos_lut[5866] = -9'sd42;
	qsin_lut[5867] =  9'sd92;
	icos_lut[5867] = -9'sd62;
	qsin_lut[5868] =  9'sd78;
	icos_lut[5868] = -9'sd78;
	qsin_lut[5869] =  9'sd62;
	icos_lut[5869] = -9'sd92;
	qsin_lut[5870] =  9'sd42;
	icos_lut[5870] = -9'sd103;
	qsin_lut[5871] =  9'sd22;
	icos_lut[5871] = -9'sd109;
	qsin_lut[5872] =  9'sd0;
	icos_lut[5872] = -9'sd111;
	qsin_lut[5873] = -9'sd22;
	icos_lut[5873] = -9'sd109;
	qsin_lut[5874] = -9'sd42;
	icos_lut[5874] = -9'sd103;
	qsin_lut[5875] = -9'sd62;
	icos_lut[5875] = -9'sd92;
	qsin_lut[5876] = -9'sd78;
	icos_lut[5876] = -9'sd78;
	qsin_lut[5877] = -9'sd92;
	icos_lut[5877] = -9'sd62;
	qsin_lut[5878] = -9'sd103;
	icos_lut[5878] = -9'sd42;
	qsin_lut[5879] = -9'sd109;
	icos_lut[5879] = -9'sd22;
	qsin_lut[5880] = -9'sd111;
	icos_lut[5880] = -9'sd0;
	qsin_lut[5881] = -9'sd109;
	icos_lut[5881] =  9'sd22;
	qsin_lut[5882] = -9'sd103;
	icos_lut[5882] =  9'sd42;
	qsin_lut[5883] = -9'sd92;
	icos_lut[5883] =  9'sd62;
	qsin_lut[5884] = -9'sd78;
	icos_lut[5884] =  9'sd78;
	qsin_lut[5885] = -9'sd62;
	icos_lut[5885] =  9'sd92;
	qsin_lut[5886] = -9'sd42;
	icos_lut[5886] =  9'sd103;
	qsin_lut[5887] = -9'sd22;
	icos_lut[5887] =  9'sd109;
	qsin_lut[5888] =  9'sd0;
	icos_lut[5888] =  9'sd113;
	qsin_lut[5889] =  9'sd22;
	icos_lut[5889] =  9'sd111;
	qsin_lut[5890] =  9'sd43;
	icos_lut[5890] =  9'sd104;
	qsin_lut[5891] =  9'sd63;
	icos_lut[5891] =  9'sd94;
	qsin_lut[5892] =  9'sd80;
	icos_lut[5892] =  9'sd80;
	qsin_lut[5893] =  9'sd94;
	icos_lut[5893] =  9'sd63;
	qsin_lut[5894] =  9'sd104;
	icos_lut[5894] =  9'sd43;
	qsin_lut[5895] =  9'sd111;
	icos_lut[5895] =  9'sd22;
	qsin_lut[5896] =  9'sd113;
	icos_lut[5896] =  9'sd0;
	qsin_lut[5897] =  9'sd111;
	icos_lut[5897] = -9'sd22;
	qsin_lut[5898] =  9'sd104;
	icos_lut[5898] = -9'sd43;
	qsin_lut[5899] =  9'sd94;
	icos_lut[5899] = -9'sd63;
	qsin_lut[5900] =  9'sd80;
	icos_lut[5900] = -9'sd80;
	qsin_lut[5901] =  9'sd63;
	icos_lut[5901] = -9'sd94;
	qsin_lut[5902] =  9'sd43;
	icos_lut[5902] = -9'sd104;
	qsin_lut[5903] =  9'sd22;
	icos_lut[5903] = -9'sd111;
	qsin_lut[5904] =  9'sd0;
	icos_lut[5904] = -9'sd113;
	qsin_lut[5905] = -9'sd22;
	icos_lut[5905] = -9'sd111;
	qsin_lut[5906] = -9'sd43;
	icos_lut[5906] = -9'sd104;
	qsin_lut[5907] = -9'sd63;
	icos_lut[5907] = -9'sd94;
	qsin_lut[5908] = -9'sd80;
	icos_lut[5908] = -9'sd80;
	qsin_lut[5909] = -9'sd94;
	icos_lut[5909] = -9'sd63;
	qsin_lut[5910] = -9'sd104;
	icos_lut[5910] = -9'sd43;
	qsin_lut[5911] = -9'sd111;
	icos_lut[5911] = -9'sd22;
	qsin_lut[5912] = -9'sd113;
	icos_lut[5912] = -9'sd0;
	qsin_lut[5913] = -9'sd111;
	icos_lut[5913] =  9'sd22;
	qsin_lut[5914] = -9'sd104;
	icos_lut[5914] =  9'sd43;
	qsin_lut[5915] = -9'sd94;
	icos_lut[5915] =  9'sd63;
	qsin_lut[5916] = -9'sd80;
	icos_lut[5916] =  9'sd80;
	qsin_lut[5917] = -9'sd63;
	icos_lut[5917] =  9'sd94;
	qsin_lut[5918] = -9'sd43;
	icos_lut[5918] =  9'sd104;
	qsin_lut[5919] = -9'sd22;
	icos_lut[5919] =  9'sd111;
	qsin_lut[5920] =  9'sd0;
	icos_lut[5920] =  9'sd115;
	qsin_lut[5921] =  9'sd22;
	icos_lut[5921] =  9'sd113;
	qsin_lut[5922] =  9'sd44;
	icos_lut[5922] =  9'sd106;
	qsin_lut[5923] =  9'sd64;
	icos_lut[5923] =  9'sd96;
	qsin_lut[5924] =  9'sd81;
	icos_lut[5924] =  9'sd81;
	qsin_lut[5925] =  9'sd96;
	icos_lut[5925] =  9'sd64;
	qsin_lut[5926] =  9'sd106;
	icos_lut[5926] =  9'sd44;
	qsin_lut[5927] =  9'sd113;
	icos_lut[5927] =  9'sd22;
	qsin_lut[5928] =  9'sd115;
	icos_lut[5928] =  9'sd0;
	qsin_lut[5929] =  9'sd113;
	icos_lut[5929] = -9'sd22;
	qsin_lut[5930] =  9'sd106;
	icos_lut[5930] = -9'sd44;
	qsin_lut[5931] =  9'sd96;
	icos_lut[5931] = -9'sd64;
	qsin_lut[5932] =  9'sd81;
	icos_lut[5932] = -9'sd81;
	qsin_lut[5933] =  9'sd64;
	icos_lut[5933] = -9'sd96;
	qsin_lut[5934] =  9'sd44;
	icos_lut[5934] = -9'sd106;
	qsin_lut[5935] =  9'sd22;
	icos_lut[5935] = -9'sd113;
	qsin_lut[5936] =  9'sd0;
	icos_lut[5936] = -9'sd115;
	qsin_lut[5937] = -9'sd22;
	icos_lut[5937] = -9'sd113;
	qsin_lut[5938] = -9'sd44;
	icos_lut[5938] = -9'sd106;
	qsin_lut[5939] = -9'sd64;
	icos_lut[5939] = -9'sd96;
	qsin_lut[5940] = -9'sd81;
	icos_lut[5940] = -9'sd81;
	qsin_lut[5941] = -9'sd96;
	icos_lut[5941] = -9'sd64;
	qsin_lut[5942] = -9'sd106;
	icos_lut[5942] = -9'sd44;
	qsin_lut[5943] = -9'sd113;
	icos_lut[5943] = -9'sd22;
	qsin_lut[5944] = -9'sd115;
	icos_lut[5944] = -9'sd0;
	qsin_lut[5945] = -9'sd113;
	icos_lut[5945] =  9'sd22;
	qsin_lut[5946] = -9'sd106;
	icos_lut[5946] =  9'sd44;
	qsin_lut[5947] = -9'sd96;
	icos_lut[5947] =  9'sd64;
	qsin_lut[5948] = -9'sd81;
	icos_lut[5948] =  9'sd81;
	qsin_lut[5949] = -9'sd64;
	icos_lut[5949] =  9'sd96;
	qsin_lut[5950] = -9'sd44;
	icos_lut[5950] =  9'sd106;
	qsin_lut[5951] = -9'sd22;
	icos_lut[5951] =  9'sd113;
	qsin_lut[5952] =  9'sd0;
	icos_lut[5952] =  9'sd117;
	qsin_lut[5953] =  9'sd23;
	icos_lut[5953] =  9'sd115;
	qsin_lut[5954] =  9'sd45;
	icos_lut[5954] =  9'sd108;
	qsin_lut[5955] =  9'sd65;
	icos_lut[5955] =  9'sd97;
	qsin_lut[5956] =  9'sd83;
	icos_lut[5956] =  9'sd83;
	qsin_lut[5957] =  9'sd97;
	icos_lut[5957] =  9'sd65;
	qsin_lut[5958] =  9'sd108;
	icos_lut[5958] =  9'sd45;
	qsin_lut[5959] =  9'sd115;
	icos_lut[5959] =  9'sd23;
	qsin_lut[5960] =  9'sd117;
	icos_lut[5960] =  9'sd0;
	qsin_lut[5961] =  9'sd115;
	icos_lut[5961] = -9'sd23;
	qsin_lut[5962] =  9'sd108;
	icos_lut[5962] = -9'sd45;
	qsin_lut[5963] =  9'sd97;
	icos_lut[5963] = -9'sd65;
	qsin_lut[5964] =  9'sd83;
	icos_lut[5964] = -9'sd83;
	qsin_lut[5965] =  9'sd65;
	icos_lut[5965] = -9'sd97;
	qsin_lut[5966] =  9'sd45;
	icos_lut[5966] = -9'sd108;
	qsin_lut[5967] =  9'sd23;
	icos_lut[5967] = -9'sd115;
	qsin_lut[5968] =  9'sd0;
	icos_lut[5968] = -9'sd117;
	qsin_lut[5969] = -9'sd23;
	icos_lut[5969] = -9'sd115;
	qsin_lut[5970] = -9'sd45;
	icos_lut[5970] = -9'sd108;
	qsin_lut[5971] = -9'sd65;
	icos_lut[5971] = -9'sd97;
	qsin_lut[5972] = -9'sd83;
	icos_lut[5972] = -9'sd83;
	qsin_lut[5973] = -9'sd97;
	icos_lut[5973] = -9'sd65;
	qsin_lut[5974] = -9'sd108;
	icos_lut[5974] = -9'sd45;
	qsin_lut[5975] = -9'sd115;
	icos_lut[5975] = -9'sd23;
	qsin_lut[5976] = -9'sd117;
	icos_lut[5976] = -9'sd0;
	qsin_lut[5977] = -9'sd115;
	icos_lut[5977] =  9'sd23;
	qsin_lut[5978] = -9'sd108;
	icos_lut[5978] =  9'sd45;
	qsin_lut[5979] = -9'sd97;
	icos_lut[5979] =  9'sd65;
	qsin_lut[5980] = -9'sd83;
	icos_lut[5980] =  9'sd83;
	qsin_lut[5981] = -9'sd65;
	icos_lut[5981] =  9'sd97;
	qsin_lut[5982] = -9'sd45;
	icos_lut[5982] =  9'sd108;
	qsin_lut[5983] = -9'sd23;
	icos_lut[5983] =  9'sd115;
	qsin_lut[5984] =  9'sd0;
	icos_lut[5984] =  9'sd119;
	qsin_lut[5985] =  9'sd23;
	icos_lut[5985] =  9'sd117;
	qsin_lut[5986] =  9'sd46;
	icos_lut[5986] =  9'sd110;
	qsin_lut[5987] =  9'sd66;
	icos_lut[5987] =  9'sd99;
	qsin_lut[5988] =  9'sd84;
	icos_lut[5988] =  9'sd84;
	qsin_lut[5989] =  9'sd99;
	icos_lut[5989] =  9'sd66;
	qsin_lut[5990] =  9'sd110;
	icos_lut[5990] =  9'sd46;
	qsin_lut[5991] =  9'sd117;
	icos_lut[5991] =  9'sd23;
	qsin_lut[5992] =  9'sd119;
	icos_lut[5992] =  9'sd0;
	qsin_lut[5993] =  9'sd117;
	icos_lut[5993] = -9'sd23;
	qsin_lut[5994] =  9'sd110;
	icos_lut[5994] = -9'sd46;
	qsin_lut[5995] =  9'sd99;
	icos_lut[5995] = -9'sd66;
	qsin_lut[5996] =  9'sd84;
	icos_lut[5996] = -9'sd84;
	qsin_lut[5997] =  9'sd66;
	icos_lut[5997] = -9'sd99;
	qsin_lut[5998] =  9'sd46;
	icos_lut[5998] = -9'sd110;
	qsin_lut[5999] =  9'sd23;
	icos_lut[5999] = -9'sd117;
	qsin_lut[6000] =  9'sd0;
	icos_lut[6000] = -9'sd119;
	qsin_lut[6001] = -9'sd23;
	icos_lut[6001] = -9'sd117;
	qsin_lut[6002] = -9'sd46;
	icos_lut[6002] = -9'sd110;
	qsin_lut[6003] = -9'sd66;
	icos_lut[6003] = -9'sd99;
	qsin_lut[6004] = -9'sd84;
	icos_lut[6004] = -9'sd84;
	qsin_lut[6005] = -9'sd99;
	icos_lut[6005] = -9'sd66;
	qsin_lut[6006] = -9'sd110;
	icos_lut[6006] = -9'sd46;
	qsin_lut[6007] = -9'sd117;
	icos_lut[6007] = -9'sd23;
	qsin_lut[6008] = -9'sd119;
	icos_lut[6008] = -9'sd0;
	qsin_lut[6009] = -9'sd117;
	icos_lut[6009] =  9'sd23;
	qsin_lut[6010] = -9'sd110;
	icos_lut[6010] =  9'sd46;
	qsin_lut[6011] = -9'sd99;
	icos_lut[6011] =  9'sd66;
	qsin_lut[6012] = -9'sd84;
	icos_lut[6012] =  9'sd84;
	qsin_lut[6013] = -9'sd66;
	icos_lut[6013] =  9'sd99;
	qsin_lut[6014] = -9'sd46;
	icos_lut[6014] =  9'sd110;
	qsin_lut[6015] = -9'sd23;
	icos_lut[6015] =  9'sd117;
	qsin_lut[6016] =  9'sd0;
	icos_lut[6016] =  9'sd121;
	qsin_lut[6017] =  9'sd24;
	icos_lut[6017] =  9'sd119;
	qsin_lut[6018] =  9'sd46;
	icos_lut[6018] =  9'sd112;
	qsin_lut[6019] =  9'sd67;
	icos_lut[6019] =  9'sd101;
	qsin_lut[6020] =  9'sd86;
	icos_lut[6020] =  9'sd86;
	qsin_lut[6021] =  9'sd101;
	icos_lut[6021] =  9'sd67;
	qsin_lut[6022] =  9'sd112;
	icos_lut[6022] =  9'sd46;
	qsin_lut[6023] =  9'sd119;
	icos_lut[6023] =  9'sd24;
	qsin_lut[6024] =  9'sd121;
	icos_lut[6024] =  9'sd0;
	qsin_lut[6025] =  9'sd119;
	icos_lut[6025] = -9'sd24;
	qsin_lut[6026] =  9'sd112;
	icos_lut[6026] = -9'sd46;
	qsin_lut[6027] =  9'sd101;
	icos_lut[6027] = -9'sd67;
	qsin_lut[6028] =  9'sd86;
	icos_lut[6028] = -9'sd86;
	qsin_lut[6029] =  9'sd67;
	icos_lut[6029] = -9'sd101;
	qsin_lut[6030] =  9'sd46;
	icos_lut[6030] = -9'sd112;
	qsin_lut[6031] =  9'sd24;
	icos_lut[6031] = -9'sd119;
	qsin_lut[6032] =  9'sd0;
	icos_lut[6032] = -9'sd121;
	qsin_lut[6033] = -9'sd24;
	icos_lut[6033] = -9'sd119;
	qsin_lut[6034] = -9'sd46;
	icos_lut[6034] = -9'sd112;
	qsin_lut[6035] = -9'sd67;
	icos_lut[6035] = -9'sd101;
	qsin_lut[6036] = -9'sd86;
	icos_lut[6036] = -9'sd86;
	qsin_lut[6037] = -9'sd101;
	icos_lut[6037] = -9'sd67;
	qsin_lut[6038] = -9'sd112;
	icos_lut[6038] = -9'sd46;
	qsin_lut[6039] = -9'sd119;
	icos_lut[6039] = -9'sd24;
	qsin_lut[6040] = -9'sd121;
	icos_lut[6040] = -9'sd0;
	qsin_lut[6041] = -9'sd119;
	icos_lut[6041] =  9'sd24;
	qsin_lut[6042] = -9'sd112;
	icos_lut[6042] =  9'sd46;
	qsin_lut[6043] = -9'sd101;
	icos_lut[6043] =  9'sd67;
	qsin_lut[6044] = -9'sd86;
	icos_lut[6044] =  9'sd86;
	qsin_lut[6045] = -9'sd67;
	icos_lut[6045] =  9'sd101;
	qsin_lut[6046] = -9'sd46;
	icos_lut[6046] =  9'sd112;
	qsin_lut[6047] = -9'sd24;
	icos_lut[6047] =  9'sd119;
	qsin_lut[6048] =  9'sd0;
	icos_lut[6048] =  9'sd123;
	qsin_lut[6049] =  9'sd24;
	icos_lut[6049] =  9'sd121;
	qsin_lut[6050] =  9'sd47;
	icos_lut[6050] =  9'sd114;
	qsin_lut[6051] =  9'sd68;
	icos_lut[6051] =  9'sd102;
	qsin_lut[6052] =  9'sd87;
	icos_lut[6052] =  9'sd87;
	qsin_lut[6053] =  9'sd102;
	icos_lut[6053] =  9'sd68;
	qsin_lut[6054] =  9'sd114;
	icos_lut[6054] =  9'sd47;
	qsin_lut[6055] =  9'sd121;
	icos_lut[6055] =  9'sd24;
	qsin_lut[6056] =  9'sd123;
	icos_lut[6056] =  9'sd0;
	qsin_lut[6057] =  9'sd121;
	icos_lut[6057] = -9'sd24;
	qsin_lut[6058] =  9'sd114;
	icos_lut[6058] = -9'sd47;
	qsin_lut[6059] =  9'sd102;
	icos_lut[6059] = -9'sd68;
	qsin_lut[6060] =  9'sd87;
	icos_lut[6060] = -9'sd87;
	qsin_lut[6061] =  9'sd68;
	icos_lut[6061] = -9'sd102;
	qsin_lut[6062] =  9'sd47;
	icos_lut[6062] = -9'sd114;
	qsin_lut[6063] =  9'sd24;
	icos_lut[6063] = -9'sd121;
	qsin_lut[6064] =  9'sd0;
	icos_lut[6064] = -9'sd123;
	qsin_lut[6065] = -9'sd24;
	icos_lut[6065] = -9'sd121;
	qsin_lut[6066] = -9'sd47;
	icos_lut[6066] = -9'sd114;
	qsin_lut[6067] = -9'sd68;
	icos_lut[6067] = -9'sd102;
	qsin_lut[6068] = -9'sd87;
	icos_lut[6068] = -9'sd87;
	qsin_lut[6069] = -9'sd102;
	icos_lut[6069] = -9'sd68;
	qsin_lut[6070] = -9'sd114;
	icos_lut[6070] = -9'sd47;
	qsin_lut[6071] = -9'sd121;
	icos_lut[6071] = -9'sd24;
	qsin_lut[6072] = -9'sd123;
	icos_lut[6072] = -9'sd0;
	qsin_lut[6073] = -9'sd121;
	icos_lut[6073] =  9'sd24;
	qsin_lut[6074] = -9'sd114;
	icos_lut[6074] =  9'sd47;
	qsin_lut[6075] = -9'sd102;
	icos_lut[6075] =  9'sd68;
	qsin_lut[6076] = -9'sd87;
	icos_lut[6076] =  9'sd87;
	qsin_lut[6077] = -9'sd68;
	icos_lut[6077] =  9'sd102;
	qsin_lut[6078] = -9'sd47;
	icos_lut[6078] =  9'sd114;
	qsin_lut[6079] = -9'sd24;
	icos_lut[6079] =  9'sd121;
	qsin_lut[6080] =  9'sd0;
	icos_lut[6080] =  9'sd125;
	qsin_lut[6081] =  9'sd24;
	icos_lut[6081] =  9'sd123;
	qsin_lut[6082] =  9'sd48;
	icos_lut[6082] =  9'sd115;
	qsin_lut[6083] =  9'sd69;
	icos_lut[6083] =  9'sd104;
	qsin_lut[6084] =  9'sd88;
	icos_lut[6084] =  9'sd88;
	qsin_lut[6085] =  9'sd104;
	icos_lut[6085] =  9'sd69;
	qsin_lut[6086] =  9'sd115;
	icos_lut[6086] =  9'sd48;
	qsin_lut[6087] =  9'sd123;
	icos_lut[6087] =  9'sd24;
	qsin_lut[6088] =  9'sd125;
	icos_lut[6088] =  9'sd0;
	qsin_lut[6089] =  9'sd123;
	icos_lut[6089] = -9'sd24;
	qsin_lut[6090] =  9'sd115;
	icos_lut[6090] = -9'sd48;
	qsin_lut[6091] =  9'sd104;
	icos_lut[6091] = -9'sd69;
	qsin_lut[6092] =  9'sd88;
	icos_lut[6092] = -9'sd88;
	qsin_lut[6093] =  9'sd69;
	icos_lut[6093] = -9'sd104;
	qsin_lut[6094] =  9'sd48;
	icos_lut[6094] = -9'sd115;
	qsin_lut[6095] =  9'sd24;
	icos_lut[6095] = -9'sd123;
	qsin_lut[6096] =  9'sd0;
	icos_lut[6096] = -9'sd125;
	qsin_lut[6097] = -9'sd24;
	icos_lut[6097] = -9'sd123;
	qsin_lut[6098] = -9'sd48;
	icos_lut[6098] = -9'sd115;
	qsin_lut[6099] = -9'sd69;
	icos_lut[6099] = -9'sd104;
	qsin_lut[6100] = -9'sd88;
	icos_lut[6100] = -9'sd88;
	qsin_lut[6101] = -9'sd104;
	icos_lut[6101] = -9'sd69;
	qsin_lut[6102] = -9'sd115;
	icos_lut[6102] = -9'sd48;
	qsin_lut[6103] = -9'sd123;
	icos_lut[6103] = -9'sd24;
	qsin_lut[6104] = -9'sd125;
	icos_lut[6104] = -9'sd0;
	qsin_lut[6105] = -9'sd123;
	icos_lut[6105] =  9'sd24;
	qsin_lut[6106] = -9'sd115;
	icos_lut[6106] =  9'sd48;
	qsin_lut[6107] = -9'sd104;
	icos_lut[6107] =  9'sd69;
	qsin_lut[6108] = -9'sd88;
	icos_lut[6108] =  9'sd88;
	qsin_lut[6109] = -9'sd69;
	icos_lut[6109] =  9'sd104;
	qsin_lut[6110] = -9'sd48;
	icos_lut[6110] =  9'sd115;
	qsin_lut[6111] = -9'sd24;
	icos_lut[6111] =  9'sd123;
	qsin_lut[6112] =  9'sd0;
	icos_lut[6112] =  9'sd127;
	qsin_lut[6113] =  9'sd25;
	icos_lut[6113] =  9'sd125;
	qsin_lut[6114] =  9'sd49;
	icos_lut[6114] =  9'sd117;
	qsin_lut[6115] =  9'sd71;
	icos_lut[6115] =  9'sd106;
	qsin_lut[6116] =  9'sd90;
	icos_lut[6116] =  9'sd90;
	qsin_lut[6117] =  9'sd106;
	icos_lut[6117] =  9'sd71;
	qsin_lut[6118] =  9'sd117;
	icos_lut[6118] =  9'sd49;
	qsin_lut[6119] =  9'sd125;
	icos_lut[6119] =  9'sd25;
	qsin_lut[6120] =  9'sd127;
	icos_lut[6120] =  9'sd0;
	qsin_lut[6121] =  9'sd125;
	icos_lut[6121] = -9'sd25;
	qsin_lut[6122] =  9'sd117;
	icos_lut[6122] = -9'sd49;
	qsin_lut[6123] =  9'sd106;
	icos_lut[6123] = -9'sd71;
	qsin_lut[6124] =  9'sd90;
	icos_lut[6124] = -9'sd90;
	qsin_lut[6125] =  9'sd71;
	icos_lut[6125] = -9'sd106;
	qsin_lut[6126] =  9'sd49;
	icos_lut[6126] = -9'sd117;
	qsin_lut[6127] =  9'sd25;
	icos_lut[6127] = -9'sd125;
	qsin_lut[6128] =  9'sd0;
	icos_lut[6128] = -9'sd127;
	qsin_lut[6129] = -9'sd25;
	icos_lut[6129] = -9'sd125;
	qsin_lut[6130] = -9'sd49;
	icos_lut[6130] = -9'sd117;
	qsin_lut[6131] = -9'sd71;
	icos_lut[6131] = -9'sd106;
	qsin_lut[6132] = -9'sd90;
	icos_lut[6132] = -9'sd90;
	qsin_lut[6133] = -9'sd106;
	icos_lut[6133] = -9'sd71;
	qsin_lut[6134] = -9'sd117;
	icos_lut[6134] = -9'sd49;
	qsin_lut[6135] = -9'sd125;
	icos_lut[6135] = -9'sd25;
	qsin_lut[6136] = -9'sd127;
	icos_lut[6136] = -9'sd0;
	qsin_lut[6137] = -9'sd125;
	icos_lut[6137] =  9'sd25;
	qsin_lut[6138] = -9'sd117;
	icos_lut[6138] =  9'sd49;
	qsin_lut[6139] = -9'sd106;
	icos_lut[6139] =  9'sd71;
	qsin_lut[6140] = -9'sd90;
	icos_lut[6140] =  9'sd90;
	qsin_lut[6141] = -9'sd71;
	icos_lut[6141] =  9'sd106;
	qsin_lut[6142] = -9'sd49;
	icos_lut[6142] =  9'sd117;
	qsin_lut[6143] = -9'sd25;
	icos_lut[6143] =  9'sd125;
	qsin_lut[6144] =  9'sd0;
	icos_lut[6144] =  9'sd129;
	qsin_lut[6145] =  9'sd25;
	icos_lut[6145] =  9'sd127;
	qsin_lut[6146] =  9'sd49;
	icos_lut[6146] =  9'sd119;
	qsin_lut[6147] =  9'sd72;
	icos_lut[6147] =  9'sd107;
	qsin_lut[6148] =  9'sd91;
	icos_lut[6148] =  9'sd91;
	qsin_lut[6149] =  9'sd107;
	icos_lut[6149] =  9'sd72;
	qsin_lut[6150] =  9'sd119;
	icos_lut[6150] =  9'sd49;
	qsin_lut[6151] =  9'sd127;
	icos_lut[6151] =  9'sd25;
	qsin_lut[6152] =  9'sd129;
	icos_lut[6152] =  9'sd0;
	qsin_lut[6153] =  9'sd127;
	icos_lut[6153] = -9'sd25;
	qsin_lut[6154] =  9'sd119;
	icos_lut[6154] = -9'sd49;
	qsin_lut[6155] =  9'sd107;
	icos_lut[6155] = -9'sd72;
	qsin_lut[6156] =  9'sd91;
	icos_lut[6156] = -9'sd91;
	qsin_lut[6157] =  9'sd72;
	icos_lut[6157] = -9'sd107;
	qsin_lut[6158] =  9'sd49;
	icos_lut[6158] = -9'sd119;
	qsin_lut[6159] =  9'sd25;
	icos_lut[6159] = -9'sd127;
	qsin_lut[6160] =  9'sd0;
	icos_lut[6160] = -9'sd129;
	qsin_lut[6161] = -9'sd25;
	icos_lut[6161] = -9'sd127;
	qsin_lut[6162] = -9'sd49;
	icos_lut[6162] = -9'sd119;
	qsin_lut[6163] = -9'sd72;
	icos_lut[6163] = -9'sd107;
	qsin_lut[6164] = -9'sd91;
	icos_lut[6164] = -9'sd91;
	qsin_lut[6165] = -9'sd107;
	icos_lut[6165] = -9'sd72;
	qsin_lut[6166] = -9'sd119;
	icos_lut[6166] = -9'sd49;
	qsin_lut[6167] = -9'sd127;
	icos_lut[6167] = -9'sd25;
	qsin_lut[6168] = -9'sd129;
	icos_lut[6168] = -9'sd0;
	qsin_lut[6169] = -9'sd127;
	icos_lut[6169] =  9'sd25;
	qsin_lut[6170] = -9'sd119;
	icos_lut[6170] =  9'sd49;
	qsin_lut[6171] = -9'sd107;
	icos_lut[6171] =  9'sd72;
	qsin_lut[6172] = -9'sd91;
	icos_lut[6172] =  9'sd91;
	qsin_lut[6173] = -9'sd72;
	icos_lut[6173] =  9'sd107;
	qsin_lut[6174] = -9'sd49;
	icos_lut[6174] =  9'sd119;
	qsin_lut[6175] = -9'sd25;
	icos_lut[6175] =  9'sd127;
	qsin_lut[6176] =  9'sd0;
	icos_lut[6176] =  9'sd131;
	qsin_lut[6177] =  9'sd26;
	icos_lut[6177] =  9'sd128;
	qsin_lut[6178] =  9'sd50;
	icos_lut[6178] =  9'sd121;
	qsin_lut[6179] =  9'sd73;
	icos_lut[6179] =  9'sd109;
	qsin_lut[6180] =  9'sd93;
	icos_lut[6180] =  9'sd93;
	qsin_lut[6181] =  9'sd109;
	icos_lut[6181] =  9'sd73;
	qsin_lut[6182] =  9'sd121;
	icos_lut[6182] =  9'sd50;
	qsin_lut[6183] =  9'sd128;
	icos_lut[6183] =  9'sd26;
	qsin_lut[6184] =  9'sd131;
	icos_lut[6184] =  9'sd0;
	qsin_lut[6185] =  9'sd128;
	icos_lut[6185] = -9'sd26;
	qsin_lut[6186] =  9'sd121;
	icos_lut[6186] = -9'sd50;
	qsin_lut[6187] =  9'sd109;
	icos_lut[6187] = -9'sd73;
	qsin_lut[6188] =  9'sd93;
	icos_lut[6188] = -9'sd93;
	qsin_lut[6189] =  9'sd73;
	icos_lut[6189] = -9'sd109;
	qsin_lut[6190] =  9'sd50;
	icos_lut[6190] = -9'sd121;
	qsin_lut[6191] =  9'sd26;
	icos_lut[6191] = -9'sd128;
	qsin_lut[6192] =  9'sd0;
	icos_lut[6192] = -9'sd131;
	qsin_lut[6193] = -9'sd26;
	icos_lut[6193] = -9'sd128;
	qsin_lut[6194] = -9'sd50;
	icos_lut[6194] = -9'sd121;
	qsin_lut[6195] = -9'sd73;
	icos_lut[6195] = -9'sd109;
	qsin_lut[6196] = -9'sd93;
	icos_lut[6196] = -9'sd93;
	qsin_lut[6197] = -9'sd109;
	icos_lut[6197] = -9'sd73;
	qsin_lut[6198] = -9'sd121;
	icos_lut[6198] = -9'sd50;
	qsin_lut[6199] = -9'sd128;
	icos_lut[6199] = -9'sd26;
	qsin_lut[6200] = -9'sd131;
	icos_lut[6200] = -9'sd0;
	qsin_lut[6201] = -9'sd128;
	icos_lut[6201] =  9'sd26;
	qsin_lut[6202] = -9'sd121;
	icos_lut[6202] =  9'sd50;
	qsin_lut[6203] = -9'sd109;
	icos_lut[6203] =  9'sd73;
	qsin_lut[6204] = -9'sd93;
	icos_lut[6204] =  9'sd93;
	qsin_lut[6205] = -9'sd73;
	icos_lut[6205] =  9'sd109;
	qsin_lut[6206] = -9'sd50;
	icos_lut[6206] =  9'sd121;
	qsin_lut[6207] = -9'sd26;
	icos_lut[6207] =  9'sd128;
	qsin_lut[6208] =  9'sd0;
	icos_lut[6208] =  9'sd133;
	qsin_lut[6209] =  9'sd26;
	icos_lut[6209] =  9'sd130;
	qsin_lut[6210] =  9'sd51;
	icos_lut[6210] =  9'sd123;
	qsin_lut[6211] =  9'sd74;
	icos_lut[6211] =  9'sd111;
	qsin_lut[6212] =  9'sd94;
	icos_lut[6212] =  9'sd94;
	qsin_lut[6213] =  9'sd111;
	icos_lut[6213] =  9'sd74;
	qsin_lut[6214] =  9'sd123;
	icos_lut[6214] =  9'sd51;
	qsin_lut[6215] =  9'sd130;
	icos_lut[6215] =  9'sd26;
	qsin_lut[6216] =  9'sd133;
	icos_lut[6216] =  9'sd0;
	qsin_lut[6217] =  9'sd130;
	icos_lut[6217] = -9'sd26;
	qsin_lut[6218] =  9'sd123;
	icos_lut[6218] = -9'sd51;
	qsin_lut[6219] =  9'sd111;
	icos_lut[6219] = -9'sd74;
	qsin_lut[6220] =  9'sd94;
	icos_lut[6220] = -9'sd94;
	qsin_lut[6221] =  9'sd74;
	icos_lut[6221] = -9'sd111;
	qsin_lut[6222] =  9'sd51;
	icos_lut[6222] = -9'sd123;
	qsin_lut[6223] =  9'sd26;
	icos_lut[6223] = -9'sd130;
	qsin_lut[6224] =  9'sd0;
	icos_lut[6224] = -9'sd133;
	qsin_lut[6225] = -9'sd26;
	icos_lut[6225] = -9'sd130;
	qsin_lut[6226] = -9'sd51;
	icos_lut[6226] = -9'sd123;
	qsin_lut[6227] = -9'sd74;
	icos_lut[6227] = -9'sd111;
	qsin_lut[6228] = -9'sd94;
	icos_lut[6228] = -9'sd94;
	qsin_lut[6229] = -9'sd111;
	icos_lut[6229] = -9'sd74;
	qsin_lut[6230] = -9'sd123;
	icos_lut[6230] = -9'sd51;
	qsin_lut[6231] = -9'sd130;
	icos_lut[6231] = -9'sd26;
	qsin_lut[6232] = -9'sd133;
	icos_lut[6232] = -9'sd0;
	qsin_lut[6233] = -9'sd130;
	icos_lut[6233] =  9'sd26;
	qsin_lut[6234] = -9'sd123;
	icos_lut[6234] =  9'sd51;
	qsin_lut[6235] = -9'sd111;
	icos_lut[6235] =  9'sd74;
	qsin_lut[6236] = -9'sd94;
	icos_lut[6236] =  9'sd94;
	qsin_lut[6237] = -9'sd74;
	icos_lut[6237] =  9'sd111;
	qsin_lut[6238] = -9'sd51;
	icos_lut[6238] =  9'sd123;
	qsin_lut[6239] = -9'sd26;
	icos_lut[6239] =  9'sd130;
	qsin_lut[6240] =  9'sd0;
	icos_lut[6240] =  9'sd135;
	qsin_lut[6241] =  9'sd26;
	icos_lut[6241] =  9'sd132;
	qsin_lut[6242] =  9'sd52;
	icos_lut[6242] =  9'sd125;
	qsin_lut[6243] =  9'sd75;
	icos_lut[6243] =  9'sd112;
	qsin_lut[6244] =  9'sd95;
	icos_lut[6244] =  9'sd95;
	qsin_lut[6245] =  9'sd112;
	icos_lut[6245] =  9'sd75;
	qsin_lut[6246] =  9'sd125;
	icos_lut[6246] =  9'sd52;
	qsin_lut[6247] =  9'sd132;
	icos_lut[6247] =  9'sd26;
	qsin_lut[6248] =  9'sd135;
	icos_lut[6248] =  9'sd0;
	qsin_lut[6249] =  9'sd132;
	icos_lut[6249] = -9'sd26;
	qsin_lut[6250] =  9'sd125;
	icos_lut[6250] = -9'sd52;
	qsin_lut[6251] =  9'sd112;
	icos_lut[6251] = -9'sd75;
	qsin_lut[6252] =  9'sd95;
	icos_lut[6252] = -9'sd95;
	qsin_lut[6253] =  9'sd75;
	icos_lut[6253] = -9'sd112;
	qsin_lut[6254] =  9'sd52;
	icos_lut[6254] = -9'sd125;
	qsin_lut[6255] =  9'sd26;
	icos_lut[6255] = -9'sd132;
	qsin_lut[6256] =  9'sd0;
	icos_lut[6256] = -9'sd135;
	qsin_lut[6257] = -9'sd26;
	icos_lut[6257] = -9'sd132;
	qsin_lut[6258] = -9'sd52;
	icos_lut[6258] = -9'sd125;
	qsin_lut[6259] = -9'sd75;
	icos_lut[6259] = -9'sd112;
	qsin_lut[6260] = -9'sd95;
	icos_lut[6260] = -9'sd95;
	qsin_lut[6261] = -9'sd112;
	icos_lut[6261] = -9'sd75;
	qsin_lut[6262] = -9'sd125;
	icos_lut[6262] = -9'sd52;
	qsin_lut[6263] = -9'sd132;
	icos_lut[6263] = -9'sd26;
	qsin_lut[6264] = -9'sd135;
	icos_lut[6264] = -9'sd0;
	qsin_lut[6265] = -9'sd132;
	icos_lut[6265] =  9'sd26;
	qsin_lut[6266] = -9'sd125;
	icos_lut[6266] =  9'sd52;
	qsin_lut[6267] = -9'sd112;
	icos_lut[6267] =  9'sd75;
	qsin_lut[6268] = -9'sd95;
	icos_lut[6268] =  9'sd95;
	qsin_lut[6269] = -9'sd75;
	icos_lut[6269] =  9'sd112;
	qsin_lut[6270] = -9'sd52;
	icos_lut[6270] =  9'sd125;
	qsin_lut[6271] = -9'sd26;
	icos_lut[6271] =  9'sd132;
	qsin_lut[6272] =  9'sd0;
	icos_lut[6272] =  9'sd137;
	qsin_lut[6273] =  9'sd27;
	icos_lut[6273] =  9'sd134;
	qsin_lut[6274] =  9'sd52;
	icos_lut[6274] =  9'sd127;
	qsin_lut[6275] =  9'sd76;
	icos_lut[6275] =  9'sd114;
	qsin_lut[6276] =  9'sd97;
	icos_lut[6276] =  9'sd97;
	qsin_lut[6277] =  9'sd114;
	icos_lut[6277] =  9'sd76;
	qsin_lut[6278] =  9'sd127;
	icos_lut[6278] =  9'sd52;
	qsin_lut[6279] =  9'sd134;
	icos_lut[6279] =  9'sd27;
	qsin_lut[6280] =  9'sd137;
	icos_lut[6280] =  9'sd0;
	qsin_lut[6281] =  9'sd134;
	icos_lut[6281] = -9'sd27;
	qsin_lut[6282] =  9'sd127;
	icos_lut[6282] = -9'sd52;
	qsin_lut[6283] =  9'sd114;
	icos_lut[6283] = -9'sd76;
	qsin_lut[6284] =  9'sd97;
	icos_lut[6284] = -9'sd97;
	qsin_lut[6285] =  9'sd76;
	icos_lut[6285] = -9'sd114;
	qsin_lut[6286] =  9'sd52;
	icos_lut[6286] = -9'sd127;
	qsin_lut[6287] =  9'sd27;
	icos_lut[6287] = -9'sd134;
	qsin_lut[6288] =  9'sd0;
	icos_lut[6288] = -9'sd137;
	qsin_lut[6289] = -9'sd27;
	icos_lut[6289] = -9'sd134;
	qsin_lut[6290] = -9'sd52;
	icos_lut[6290] = -9'sd127;
	qsin_lut[6291] = -9'sd76;
	icos_lut[6291] = -9'sd114;
	qsin_lut[6292] = -9'sd97;
	icos_lut[6292] = -9'sd97;
	qsin_lut[6293] = -9'sd114;
	icos_lut[6293] = -9'sd76;
	qsin_lut[6294] = -9'sd127;
	icos_lut[6294] = -9'sd52;
	qsin_lut[6295] = -9'sd134;
	icos_lut[6295] = -9'sd27;
	qsin_lut[6296] = -9'sd137;
	icos_lut[6296] = -9'sd0;
	qsin_lut[6297] = -9'sd134;
	icos_lut[6297] =  9'sd27;
	qsin_lut[6298] = -9'sd127;
	icos_lut[6298] =  9'sd52;
	qsin_lut[6299] = -9'sd114;
	icos_lut[6299] =  9'sd76;
	qsin_lut[6300] = -9'sd97;
	icos_lut[6300] =  9'sd97;
	qsin_lut[6301] = -9'sd76;
	icos_lut[6301] =  9'sd114;
	qsin_lut[6302] = -9'sd52;
	icos_lut[6302] =  9'sd127;
	qsin_lut[6303] = -9'sd27;
	icos_lut[6303] =  9'sd134;
	qsin_lut[6304] =  9'sd0;
	icos_lut[6304] =  9'sd139;
	qsin_lut[6305] =  9'sd27;
	icos_lut[6305] =  9'sd136;
	qsin_lut[6306] =  9'sd53;
	icos_lut[6306] =  9'sd128;
	qsin_lut[6307] =  9'sd77;
	icos_lut[6307] =  9'sd116;
	qsin_lut[6308] =  9'sd98;
	icos_lut[6308] =  9'sd98;
	qsin_lut[6309] =  9'sd116;
	icos_lut[6309] =  9'sd77;
	qsin_lut[6310] =  9'sd128;
	icos_lut[6310] =  9'sd53;
	qsin_lut[6311] =  9'sd136;
	icos_lut[6311] =  9'sd27;
	qsin_lut[6312] =  9'sd139;
	icos_lut[6312] =  9'sd0;
	qsin_lut[6313] =  9'sd136;
	icos_lut[6313] = -9'sd27;
	qsin_lut[6314] =  9'sd128;
	icos_lut[6314] = -9'sd53;
	qsin_lut[6315] =  9'sd116;
	icos_lut[6315] = -9'sd77;
	qsin_lut[6316] =  9'sd98;
	icos_lut[6316] = -9'sd98;
	qsin_lut[6317] =  9'sd77;
	icos_lut[6317] = -9'sd116;
	qsin_lut[6318] =  9'sd53;
	icos_lut[6318] = -9'sd128;
	qsin_lut[6319] =  9'sd27;
	icos_lut[6319] = -9'sd136;
	qsin_lut[6320] =  9'sd0;
	icos_lut[6320] = -9'sd139;
	qsin_lut[6321] = -9'sd27;
	icos_lut[6321] = -9'sd136;
	qsin_lut[6322] = -9'sd53;
	icos_lut[6322] = -9'sd128;
	qsin_lut[6323] = -9'sd77;
	icos_lut[6323] = -9'sd116;
	qsin_lut[6324] = -9'sd98;
	icos_lut[6324] = -9'sd98;
	qsin_lut[6325] = -9'sd116;
	icos_lut[6325] = -9'sd77;
	qsin_lut[6326] = -9'sd128;
	icos_lut[6326] = -9'sd53;
	qsin_lut[6327] = -9'sd136;
	icos_lut[6327] = -9'sd27;
	qsin_lut[6328] = -9'sd139;
	icos_lut[6328] = -9'sd0;
	qsin_lut[6329] = -9'sd136;
	icos_lut[6329] =  9'sd27;
	qsin_lut[6330] = -9'sd128;
	icos_lut[6330] =  9'sd53;
	qsin_lut[6331] = -9'sd116;
	icos_lut[6331] =  9'sd77;
	qsin_lut[6332] = -9'sd98;
	icos_lut[6332] =  9'sd98;
	qsin_lut[6333] = -9'sd77;
	icos_lut[6333] =  9'sd116;
	qsin_lut[6334] = -9'sd53;
	icos_lut[6334] =  9'sd128;
	qsin_lut[6335] = -9'sd27;
	icos_lut[6335] =  9'sd136;
	qsin_lut[6336] =  9'sd0;
	icos_lut[6336] =  9'sd141;
	qsin_lut[6337] =  9'sd28;
	icos_lut[6337] =  9'sd138;
	qsin_lut[6338] =  9'sd54;
	icos_lut[6338] =  9'sd130;
	qsin_lut[6339] =  9'sd78;
	icos_lut[6339] =  9'sd117;
	qsin_lut[6340] =  9'sd100;
	icos_lut[6340] =  9'sd100;
	qsin_lut[6341] =  9'sd117;
	icos_lut[6341] =  9'sd78;
	qsin_lut[6342] =  9'sd130;
	icos_lut[6342] =  9'sd54;
	qsin_lut[6343] =  9'sd138;
	icos_lut[6343] =  9'sd28;
	qsin_lut[6344] =  9'sd141;
	icos_lut[6344] =  9'sd0;
	qsin_lut[6345] =  9'sd138;
	icos_lut[6345] = -9'sd28;
	qsin_lut[6346] =  9'sd130;
	icos_lut[6346] = -9'sd54;
	qsin_lut[6347] =  9'sd117;
	icos_lut[6347] = -9'sd78;
	qsin_lut[6348] =  9'sd100;
	icos_lut[6348] = -9'sd100;
	qsin_lut[6349] =  9'sd78;
	icos_lut[6349] = -9'sd117;
	qsin_lut[6350] =  9'sd54;
	icos_lut[6350] = -9'sd130;
	qsin_lut[6351] =  9'sd28;
	icos_lut[6351] = -9'sd138;
	qsin_lut[6352] =  9'sd0;
	icos_lut[6352] = -9'sd141;
	qsin_lut[6353] = -9'sd28;
	icos_lut[6353] = -9'sd138;
	qsin_lut[6354] = -9'sd54;
	icos_lut[6354] = -9'sd130;
	qsin_lut[6355] = -9'sd78;
	icos_lut[6355] = -9'sd117;
	qsin_lut[6356] = -9'sd100;
	icos_lut[6356] = -9'sd100;
	qsin_lut[6357] = -9'sd117;
	icos_lut[6357] = -9'sd78;
	qsin_lut[6358] = -9'sd130;
	icos_lut[6358] = -9'sd54;
	qsin_lut[6359] = -9'sd138;
	icos_lut[6359] = -9'sd28;
	qsin_lut[6360] = -9'sd141;
	icos_lut[6360] = -9'sd0;
	qsin_lut[6361] = -9'sd138;
	icos_lut[6361] =  9'sd28;
	qsin_lut[6362] = -9'sd130;
	icos_lut[6362] =  9'sd54;
	qsin_lut[6363] = -9'sd117;
	icos_lut[6363] =  9'sd78;
	qsin_lut[6364] = -9'sd100;
	icos_lut[6364] =  9'sd100;
	qsin_lut[6365] = -9'sd78;
	icos_lut[6365] =  9'sd117;
	qsin_lut[6366] = -9'sd54;
	icos_lut[6366] =  9'sd130;
	qsin_lut[6367] = -9'sd28;
	icos_lut[6367] =  9'sd138;
	qsin_lut[6368] =  9'sd0;
	icos_lut[6368] =  9'sd143;
	qsin_lut[6369] =  9'sd28;
	icos_lut[6369] =  9'sd140;
	qsin_lut[6370] =  9'sd55;
	icos_lut[6370] =  9'sd132;
	qsin_lut[6371] =  9'sd79;
	icos_lut[6371] =  9'sd119;
	qsin_lut[6372] =  9'sd101;
	icos_lut[6372] =  9'sd101;
	qsin_lut[6373] =  9'sd119;
	icos_lut[6373] =  9'sd79;
	qsin_lut[6374] =  9'sd132;
	icos_lut[6374] =  9'sd55;
	qsin_lut[6375] =  9'sd140;
	icos_lut[6375] =  9'sd28;
	qsin_lut[6376] =  9'sd143;
	icos_lut[6376] =  9'sd0;
	qsin_lut[6377] =  9'sd140;
	icos_lut[6377] = -9'sd28;
	qsin_lut[6378] =  9'sd132;
	icos_lut[6378] = -9'sd55;
	qsin_lut[6379] =  9'sd119;
	icos_lut[6379] = -9'sd79;
	qsin_lut[6380] =  9'sd101;
	icos_lut[6380] = -9'sd101;
	qsin_lut[6381] =  9'sd79;
	icos_lut[6381] = -9'sd119;
	qsin_lut[6382] =  9'sd55;
	icos_lut[6382] = -9'sd132;
	qsin_lut[6383] =  9'sd28;
	icos_lut[6383] = -9'sd140;
	qsin_lut[6384] =  9'sd0;
	icos_lut[6384] = -9'sd143;
	qsin_lut[6385] = -9'sd28;
	icos_lut[6385] = -9'sd140;
	qsin_lut[6386] = -9'sd55;
	icos_lut[6386] = -9'sd132;
	qsin_lut[6387] = -9'sd79;
	icos_lut[6387] = -9'sd119;
	qsin_lut[6388] = -9'sd101;
	icos_lut[6388] = -9'sd101;
	qsin_lut[6389] = -9'sd119;
	icos_lut[6389] = -9'sd79;
	qsin_lut[6390] = -9'sd132;
	icos_lut[6390] = -9'sd55;
	qsin_lut[6391] = -9'sd140;
	icos_lut[6391] = -9'sd28;
	qsin_lut[6392] = -9'sd143;
	icos_lut[6392] = -9'sd0;
	qsin_lut[6393] = -9'sd140;
	icos_lut[6393] =  9'sd28;
	qsin_lut[6394] = -9'sd132;
	icos_lut[6394] =  9'sd55;
	qsin_lut[6395] = -9'sd119;
	icos_lut[6395] =  9'sd79;
	qsin_lut[6396] = -9'sd101;
	icos_lut[6396] =  9'sd101;
	qsin_lut[6397] = -9'sd79;
	icos_lut[6397] =  9'sd119;
	qsin_lut[6398] = -9'sd55;
	icos_lut[6398] =  9'sd132;
	qsin_lut[6399] = -9'sd28;
	icos_lut[6399] =  9'sd140;
	qsin_lut[6400] =  9'sd0;
	icos_lut[6400] =  9'sd145;
	qsin_lut[6401] =  9'sd28;
	icos_lut[6401] =  9'sd142;
	qsin_lut[6402] =  9'sd55;
	icos_lut[6402] =  9'sd134;
	qsin_lut[6403] =  9'sd81;
	icos_lut[6403] =  9'sd121;
	qsin_lut[6404] =  9'sd103;
	icos_lut[6404] =  9'sd103;
	qsin_lut[6405] =  9'sd121;
	icos_lut[6405] =  9'sd81;
	qsin_lut[6406] =  9'sd134;
	icos_lut[6406] =  9'sd55;
	qsin_lut[6407] =  9'sd142;
	icos_lut[6407] =  9'sd28;
	qsin_lut[6408] =  9'sd145;
	icos_lut[6408] =  9'sd0;
	qsin_lut[6409] =  9'sd142;
	icos_lut[6409] = -9'sd28;
	qsin_lut[6410] =  9'sd134;
	icos_lut[6410] = -9'sd55;
	qsin_lut[6411] =  9'sd121;
	icos_lut[6411] = -9'sd81;
	qsin_lut[6412] =  9'sd103;
	icos_lut[6412] = -9'sd103;
	qsin_lut[6413] =  9'sd81;
	icos_lut[6413] = -9'sd121;
	qsin_lut[6414] =  9'sd55;
	icos_lut[6414] = -9'sd134;
	qsin_lut[6415] =  9'sd28;
	icos_lut[6415] = -9'sd142;
	qsin_lut[6416] =  9'sd0;
	icos_lut[6416] = -9'sd145;
	qsin_lut[6417] = -9'sd28;
	icos_lut[6417] = -9'sd142;
	qsin_lut[6418] = -9'sd55;
	icos_lut[6418] = -9'sd134;
	qsin_lut[6419] = -9'sd81;
	icos_lut[6419] = -9'sd121;
	qsin_lut[6420] = -9'sd103;
	icos_lut[6420] = -9'sd103;
	qsin_lut[6421] = -9'sd121;
	icos_lut[6421] = -9'sd81;
	qsin_lut[6422] = -9'sd134;
	icos_lut[6422] = -9'sd55;
	qsin_lut[6423] = -9'sd142;
	icos_lut[6423] = -9'sd28;
	qsin_lut[6424] = -9'sd145;
	icos_lut[6424] = -9'sd0;
	qsin_lut[6425] = -9'sd142;
	icos_lut[6425] =  9'sd28;
	qsin_lut[6426] = -9'sd134;
	icos_lut[6426] =  9'sd55;
	qsin_lut[6427] = -9'sd121;
	icos_lut[6427] =  9'sd81;
	qsin_lut[6428] = -9'sd103;
	icos_lut[6428] =  9'sd103;
	qsin_lut[6429] = -9'sd81;
	icos_lut[6429] =  9'sd121;
	qsin_lut[6430] = -9'sd55;
	icos_lut[6430] =  9'sd134;
	qsin_lut[6431] = -9'sd28;
	icos_lut[6431] =  9'sd142;
	qsin_lut[6432] =  9'sd0;
	icos_lut[6432] =  9'sd147;
	qsin_lut[6433] =  9'sd29;
	icos_lut[6433] =  9'sd144;
	qsin_lut[6434] =  9'sd56;
	icos_lut[6434] =  9'sd136;
	qsin_lut[6435] =  9'sd82;
	icos_lut[6435] =  9'sd122;
	qsin_lut[6436] =  9'sd104;
	icos_lut[6436] =  9'sd104;
	qsin_lut[6437] =  9'sd122;
	icos_lut[6437] =  9'sd82;
	qsin_lut[6438] =  9'sd136;
	icos_lut[6438] =  9'sd56;
	qsin_lut[6439] =  9'sd144;
	icos_lut[6439] =  9'sd29;
	qsin_lut[6440] =  9'sd147;
	icos_lut[6440] =  9'sd0;
	qsin_lut[6441] =  9'sd144;
	icos_lut[6441] = -9'sd29;
	qsin_lut[6442] =  9'sd136;
	icos_lut[6442] = -9'sd56;
	qsin_lut[6443] =  9'sd122;
	icos_lut[6443] = -9'sd82;
	qsin_lut[6444] =  9'sd104;
	icos_lut[6444] = -9'sd104;
	qsin_lut[6445] =  9'sd82;
	icos_lut[6445] = -9'sd122;
	qsin_lut[6446] =  9'sd56;
	icos_lut[6446] = -9'sd136;
	qsin_lut[6447] =  9'sd29;
	icos_lut[6447] = -9'sd144;
	qsin_lut[6448] =  9'sd0;
	icos_lut[6448] = -9'sd147;
	qsin_lut[6449] = -9'sd29;
	icos_lut[6449] = -9'sd144;
	qsin_lut[6450] = -9'sd56;
	icos_lut[6450] = -9'sd136;
	qsin_lut[6451] = -9'sd82;
	icos_lut[6451] = -9'sd122;
	qsin_lut[6452] = -9'sd104;
	icos_lut[6452] = -9'sd104;
	qsin_lut[6453] = -9'sd122;
	icos_lut[6453] = -9'sd82;
	qsin_lut[6454] = -9'sd136;
	icos_lut[6454] = -9'sd56;
	qsin_lut[6455] = -9'sd144;
	icos_lut[6455] = -9'sd29;
	qsin_lut[6456] = -9'sd147;
	icos_lut[6456] = -9'sd0;
	qsin_lut[6457] = -9'sd144;
	icos_lut[6457] =  9'sd29;
	qsin_lut[6458] = -9'sd136;
	icos_lut[6458] =  9'sd56;
	qsin_lut[6459] = -9'sd122;
	icos_lut[6459] =  9'sd82;
	qsin_lut[6460] = -9'sd104;
	icos_lut[6460] =  9'sd104;
	qsin_lut[6461] = -9'sd82;
	icos_lut[6461] =  9'sd122;
	qsin_lut[6462] = -9'sd56;
	icos_lut[6462] =  9'sd136;
	qsin_lut[6463] = -9'sd29;
	icos_lut[6463] =  9'sd144;
	qsin_lut[6464] =  9'sd0;
	icos_lut[6464] =  9'sd149;
	qsin_lut[6465] =  9'sd29;
	icos_lut[6465] =  9'sd146;
	qsin_lut[6466] =  9'sd57;
	icos_lut[6466] =  9'sd138;
	qsin_lut[6467] =  9'sd83;
	icos_lut[6467] =  9'sd124;
	qsin_lut[6468] =  9'sd105;
	icos_lut[6468] =  9'sd105;
	qsin_lut[6469] =  9'sd124;
	icos_lut[6469] =  9'sd83;
	qsin_lut[6470] =  9'sd138;
	icos_lut[6470] =  9'sd57;
	qsin_lut[6471] =  9'sd146;
	icos_lut[6471] =  9'sd29;
	qsin_lut[6472] =  9'sd149;
	icos_lut[6472] =  9'sd0;
	qsin_lut[6473] =  9'sd146;
	icos_lut[6473] = -9'sd29;
	qsin_lut[6474] =  9'sd138;
	icos_lut[6474] = -9'sd57;
	qsin_lut[6475] =  9'sd124;
	icos_lut[6475] = -9'sd83;
	qsin_lut[6476] =  9'sd105;
	icos_lut[6476] = -9'sd105;
	qsin_lut[6477] =  9'sd83;
	icos_lut[6477] = -9'sd124;
	qsin_lut[6478] =  9'sd57;
	icos_lut[6478] = -9'sd138;
	qsin_lut[6479] =  9'sd29;
	icos_lut[6479] = -9'sd146;
	qsin_lut[6480] =  9'sd0;
	icos_lut[6480] = -9'sd149;
	qsin_lut[6481] = -9'sd29;
	icos_lut[6481] = -9'sd146;
	qsin_lut[6482] = -9'sd57;
	icos_lut[6482] = -9'sd138;
	qsin_lut[6483] = -9'sd83;
	icos_lut[6483] = -9'sd124;
	qsin_lut[6484] = -9'sd105;
	icos_lut[6484] = -9'sd105;
	qsin_lut[6485] = -9'sd124;
	icos_lut[6485] = -9'sd83;
	qsin_lut[6486] = -9'sd138;
	icos_lut[6486] = -9'sd57;
	qsin_lut[6487] = -9'sd146;
	icos_lut[6487] = -9'sd29;
	qsin_lut[6488] = -9'sd149;
	icos_lut[6488] = -9'sd0;
	qsin_lut[6489] = -9'sd146;
	icos_lut[6489] =  9'sd29;
	qsin_lut[6490] = -9'sd138;
	icos_lut[6490] =  9'sd57;
	qsin_lut[6491] = -9'sd124;
	icos_lut[6491] =  9'sd83;
	qsin_lut[6492] = -9'sd105;
	icos_lut[6492] =  9'sd105;
	qsin_lut[6493] = -9'sd83;
	icos_lut[6493] =  9'sd124;
	qsin_lut[6494] = -9'sd57;
	icos_lut[6494] =  9'sd138;
	qsin_lut[6495] = -9'sd29;
	icos_lut[6495] =  9'sd146;
	qsin_lut[6496] =  9'sd0;
	icos_lut[6496] =  9'sd151;
	qsin_lut[6497] =  9'sd29;
	icos_lut[6497] =  9'sd148;
	qsin_lut[6498] =  9'sd58;
	icos_lut[6498] =  9'sd140;
	qsin_lut[6499] =  9'sd84;
	icos_lut[6499] =  9'sd126;
	qsin_lut[6500] =  9'sd107;
	icos_lut[6500] =  9'sd107;
	qsin_lut[6501] =  9'sd126;
	icos_lut[6501] =  9'sd84;
	qsin_lut[6502] =  9'sd140;
	icos_lut[6502] =  9'sd58;
	qsin_lut[6503] =  9'sd148;
	icos_lut[6503] =  9'sd29;
	qsin_lut[6504] =  9'sd151;
	icos_lut[6504] =  9'sd0;
	qsin_lut[6505] =  9'sd148;
	icos_lut[6505] = -9'sd29;
	qsin_lut[6506] =  9'sd140;
	icos_lut[6506] = -9'sd58;
	qsin_lut[6507] =  9'sd126;
	icos_lut[6507] = -9'sd84;
	qsin_lut[6508] =  9'sd107;
	icos_lut[6508] = -9'sd107;
	qsin_lut[6509] =  9'sd84;
	icos_lut[6509] = -9'sd126;
	qsin_lut[6510] =  9'sd58;
	icos_lut[6510] = -9'sd140;
	qsin_lut[6511] =  9'sd29;
	icos_lut[6511] = -9'sd148;
	qsin_lut[6512] =  9'sd0;
	icos_lut[6512] = -9'sd151;
	qsin_lut[6513] = -9'sd29;
	icos_lut[6513] = -9'sd148;
	qsin_lut[6514] = -9'sd58;
	icos_lut[6514] = -9'sd140;
	qsin_lut[6515] = -9'sd84;
	icos_lut[6515] = -9'sd126;
	qsin_lut[6516] = -9'sd107;
	icos_lut[6516] = -9'sd107;
	qsin_lut[6517] = -9'sd126;
	icos_lut[6517] = -9'sd84;
	qsin_lut[6518] = -9'sd140;
	icos_lut[6518] = -9'sd58;
	qsin_lut[6519] = -9'sd148;
	icos_lut[6519] = -9'sd29;
	qsin_lut[6520] = -9'sd151;
	icos_lut[6520] = -9'sd0;
	qsin_lut[6521] = -9'sd148;
	icos_lut[6521] =  9'sd29;
	qsin_lut[6522] = -9'sd140;
	icos_lut[6522] =  9'sd58;
	qsin_lut[6523] = -9'sd126;
	icos_lut[6523] =  9'sd84;
	qsin_lut[6524] = -9'sd107;
	icos_lut[6524] =  9'sd107;
	qsin_lut[6525] = -9'sd84;
	icos_lut[6525] =  9'sd126;
	qsin_lut[6526] = -9'sd58;
	icos_lut[6526] =  9'sd140;
	qsin_lut[6527] = -9'sd29;
	icos_lut[6527] =  9'sd148;
	qsin_lut[6528] =  9'sd0;
	icos_lut[6528] =  9'sd153;
	qsin_lut[6529] =  9'sd30;
	icos_lut[6529] =  9'sd150;
	qsin_lut[6530] =  9'sd59;
	icos_lut[6530] =  9'sd141;
	qsin_lut[6531] =  9'sd85;
	icos_lut[6531] =  9'sd127;
	qsin_lut[6532] =  9'sd108;
	icos_lut[6532] =  9'sd108;
	qsin_lut[6533] =  9'sd127;
	icos_lut[6533] =  9'sd85;
	qsin_lut[6534] =  9'sd141;
	icos_lut[6534] =  9'sd59;
	qsin_lut[6535] =  9'sd150;
	icos_lut[6535] =  9'sd30;
	qsin_lut[6536] =  9'sd153;
	icos_lut[6536] =  9'sd0;
	qsin_lut[6537] =  9'sd150;
	icos_lut[6537] = -9'sd30;
	qsin_lut[6538] =  9'sd141;
	icos_lut[6538] = -9'sd59;
	qsin_lut[6539] =  9'sd127;
	icos_lut[6539] = -9'sd85;
	qsin_lut[6540] =  9'sd108;
	icos_lut[6540] = -9'sd108;
	qsin_lut[6541] =  9'sd85;
	icos_lut[6541] = -9'sd127;
	qsin_lut[6542] =  9'sd59;
	icos_lut[6542] = -9'sd141;
	qsin_lut[6543] =  9'sd30;
	icos_lut[6543] = -9'sd150;
	qsin_lut[6544] =  9'sd0;
	icos_lut[6544] = -9'sd153;
	qsin_lut[6545] = -9'sd30;
	icos_lut[6545] = -9'sd150;
	qsin_lut[6546] = -9'sd59;
	icos_lut[6546] = -9'sd141;
	qsin_lut[6547] = -9'sd85;
	icos_lut[6547] = -9'sd127;
	qsin_lut[6548] = -9'sd108;
	icos_lut[6548] = -9'sd108;
	qsin_lut[6549] = -9'sd127;
	icos_lut[6549] = -9'sd85;
	qsin_lut[6550] = -9'sd141;
	icos_lut[6550] = -9'sd59;
	qsin_lut[6551] = -9'sd150;
	icos_lut[6551] = -9'sd30;
	qsin_lut[6552] = -9'sd153;
	icos_lut[6552] = -9'sd0;
	qsin_lut[6553] = -9'sd150;
	icos_lut[6553] =  9'sd30;
	qsin_lut[6554] = -9'sd141;
	icos_lut[6554] =  9'sd59;
	qsin_lut[6555] = -9'sd127;
	icos_lut[6555] =  9'sd85;
	qsin_lut[6556] = -9'sd108;
	icos_lut[6556] =  9'sd108;
	qsin_lut[6557] = -9'sd85;
	icos_lut[6557] =  9'sd127;
	qsin_lut[6558] = -9'sd59;
	icos_lut[6558] =  9'sd141;
	qsin_lut[6559] = -9'sd30;
	icos_lut[6559] =  9'sd150;
	qsin_lut[6560] =  9'sd0;
	icos_lut[6560] =  9'sd155;
	qsin_lut[6561] =  9'sd30;
	icos_lut[6561] =  9'sd152;
	qsin_lut[6562] =  9'sd59;
	icos_lut[6562] =  9'sd143;
	qsin_lut[6563] =  9'sd86;
	icos_lut[6563] =  9'sd129;
	qsin_lut[6564] =  9'sd110;
	icos_lut[6564] =  9'sd110;
	qsin_lut[6565] =  9'sd129;
	icos_lut[6565] =  9'sd86;
	qsin_lut[6566] =  9'sd143;
	icos_lut[6566] =  9'sd59;
	qsin_lut[6567] =  9'sd152;
	icos_lut[6567] =  9'sd30;
	qsin_lut[6568] =  9'sd155;
	icos_lut[6568] =  9'sd0;
	qsin_lut[6569] =  9'sd152;
	icos_lut[6569] = -9'sd30;
	qsin_lut[6570] =  9'sd143;
	icos_lut[6570] = -9'sd59;
	qsin_lut[6571] =  9'sd129;
	icos_lut[6571] = -9'sd86;
	qsin_lut[6572] =  9'sd110;
	icos_lut[6572] = -9'sd110;
	qsin_lut[6573] =  9'sd86;
	icos_lut[6573] = -9'sd129;
	qsin_lut[6574] =  9'sd59;
	icos_lut[6574] = -9'sd143;
	qsin_lut[6575] =  9'sd30;
	icos_lut[6575] = -9'sd152;
	qsin_lut[6576] =  9'sd0;
	icos_lut[6576] = -9'sd155;
	qsin_lut[6577] = -9'sd30;
	icos_lut[6577] = -9'sd152;
	qsin_lut[6578] = -9'sd59;
	icos_lut[6578] = -9'sd143;
	qsin_lut[6579] = -9'sd86;
	icos_lut[6579] = -9'sd129;
	qsin_lut[6580] = -9'sd110;
	icos_lut[6580] = -9'sd110;
	qsin_lut[6581] = -9'sd129;
	icos_lut[6581] = -9'sd86;
	qsin_lut[6582] = -9'sd143;
	icos_lut[6582] = -9'sd59;
	qsin_lut[6583] = -9'sd152;
	icos_lut[6583] = -9'sd30;
	qsin_lut[6584] = -9'sd155;
	icos_lut[6584] = -9'sd0;
	qsin_lut[6585] = -9'sd152;
	icos_lut[6585] =  9'sd30;
	qsin_lut[6586] = -9'sd143;
	icos_lut[6586] =  9'sd59;
	qsin_lut[6587] = -9'sd129;
	icos_lut[6587] =  9'sd86;
	qsin_lut[6588] = -9'sd110;
	icos_lut[6588] =  9'sd110;
	qsin_lut[6589] = -9'sd86;
	icos_lut[6589] =  9'sd129;
	qsin_lut[6590] = -9'sd59;
	icos_lut[6590] =  9'sd143;
	qsin_lut[6591] = -9'sd30;
	icos_lut[6591] =  9'sd152;
	qsin_lut[6592] =  9'sd0;
	icos_lut[6592] =  9'sd157;
	qsin_lut[6593] =  9'sd31;
	icos_lut[6593] =  9'sd154;
	qsin_lut[6594] =  9'sd60;
	icos_lut[6594] =  9'sd145;
	qsin_lut[6595] =  9'sd87;
	icos_lut[6595] =  9'sd131;
	qsin_lut[6596] =  9'sd111;
	icos_lut[6596] =  9'sd111;
	qsin_lut[6597] =  9'sd131;
	icos_lut[6597] =  9'sd87;
	qsin_lut[6598] =  9'sd145;
	icos_lut[6598] =  9'sd60;
	qsin_lut[6599] =  9'sd154;
	icos_lut[6599] =  9'sd31;
	qsin_lut[6600] =  9'sd157;
	icos_lut[6600] =  9'sd0;
	qsin_lut[6601] =  9'sd154;
	icos_lut[6601] = -9'sd31;
	qsin_lut[6602] =  9'sd145;
	icos_lut[6602] = -9'sd60;
	qsin_lut[6603] =  9'sd131;
	icos_lut[6603] = -9'sd87;
	qsin_lut[6604] =  9'sd111;
	icos_lut[6604] = -9'sd111;
	qsin_lut[6605] =  9'sd87;
	icos_lut[6605] = -9'sd131;
	qsin_lut[6606] =  9'sd60;
	icos_lut[6606] = -9'sd145;
	qsin_lut[6607] =  9'sd31;
	icos_lut[6607] = -9'sd154;
	qsin_lut[6608] =  9'sd0;
	icos_lut[6608] = -9'sd157;
	qsin_lut[6609] = -9'sd31;
	icos_lut[6609] = -9'sd154;
	qsin_lut[6610] = -9'sd60;
	icos_lut[6610] = -9'sd145;
	qsin_lut[6611] = -9'sd87;
	icos_lut[6611] = -9'sd131;
	qsin_lut[6612] = -9'sd111;
	icos_lut[6612] = -9'sd111;
	qsin_lut[6613] = -9'sd131;
	icos_lut[6613] = -9'sd87;
	qsin_lut[6614] = -9'sd145;
	icos_lut[6614] = -9'sd60;
	qsin_lut[6615] = -9'sd154;
	icos_lut[6615] = -9'sd31;
	qsin_lut[6616] = -9'sd157;
	icos_lut[6616] = -9'sd0;
	qsin_lut[6617] = -9'sd154;
	icos_lut[6617] =  9'sd31;
	qsin_lut[6618] = -9'sd145;
	icos_lut[6618] =  9'sd60;
	qsin_lut[6619] = -9'sd131;
	icos_lut[6619] =  9'sd87;
	qsin_lut[6620] = -9'sd111;
	icos_lut[6620] =  9'sd111;
	qsin_lut[6621] = -9'sd87;
	icos_lut[6621] =  9'sd131;
	qsin_lut[6622] = -9'sd60;
	icos_lut[6622] =  9'sd145;
	qsin_lut[6623] = -9'sd31;
	icos_lut[6623] =  9'sd154;
	qsin_lut[6624] =  9'sd0;
	icos_lut[6624] =  9'sd159;
	qsin_lut[6625] =  9'sd31;
	icos_lut[6625] =  9'sd156;
	qsin_lut[6626] =  9'sd61;
	icos_lut[6626] =  9'sd147;
	qsin_lut[6627] =  9'sd88;
	icos_lut[6627] =  9'sd132;
	qsin_lut[6628] =  9'sd112;
	icos_lut[6628] =  9'sd112;
	qsin_lut[6629] =  9'sd132;
	icos_lut[6629] =  9'sd88;
	qsin_lut[6630] =  9'sd147;
	icos_lut[6630] =  9'sd61;
	qsin_lut[6631] =  9'sd156;
	icos_lut[6631] =  9'sd31;
	qsin_lut[6632] =  9'sd159;
	icos_lut[6632] =  9'sd0;
	qsin_lut[6633] =  9'sd156;
	icos_lut[6633] = -9'sd31;
	qsin_lut[6634] =  9'sd147;
	icos_lut[6634] = -9'sd61;
	qsin_lut[6635] =  9'sd132;
	icos_lut[6635] = -9'sd88;
	qsin_lut[6636] =  9'sd112;
	icos_lut[6636] = -9'sd112;
	qsin_lut[6637] =  9'sd88;
	icos_lut[6637] = -9'sd132;
	qsin_lut[6638] =  9'sd61;
	icos_lut[6638] = -9'sd147;
	qsin_lut[6639] =  9'sd31;
	icos_lut[6639] = -9'sd156;
	qsin_lut[6640] =  9'sd0;
	icos_lut[6640] = -9'sd159;
	qsin_lut[6641] = -9'sd31;
	icos_lut[6641] = -9'sd156;
	qsin_lut[6642] = -9'sd61;
	icos_lut[6642] = -9'sd147;
	qsin_lut[6643] = -9'sd88;
	icos_lut[6643] = -9'sd132;
	qsin_lut[6644] = -9'sd112;
	icos_lut[6644] = -9'sd112;
	qsin_lut[6645] = -9'sd132;
	icos_lut[6645] = -9'sd88;
	qsin_lut[6646] = -9'sd147;
	icos_lut[6646] = -9'sd61;
	qsin_lut[6647] = -9'sd156;
	icos_lut[6647] = -9'sd31;
	qsin_lut[6648] = -9'sd159;
	icos_lut[6648] = -9'sd0;
	qsin_lut[6649] = -9'sd156;
	icos_lut[6649] =  9'sd31;
	qsin_lut[6650] = -9'sd147;
	icos_lut[6650] =  9'sd61;
	qsin_lut[6651] = -9'sd132;
	icos_lut[6651] =  9'sd88;
	qsin_lut[6652] = -9'sd112;
	icos_lut[6652] =  9'sd112;
	qsin_lut[6653] = -9'sd88;
	icos_lut[6653] =  9'sd132;
	qsin_lut[6654] = -9'sd61;
	icos_lut[6654] =  9'sd147;
	qsin_lut[6655] = -9'sd31;
	icos_lut[6655] =  9'sd156;
	qsin_lut[6656] =  9'sd0;
	icos_lut[6656] =  9'sd161;
	qsin_lut[6657] =  9'sd31;
	icos_lut[6657] =  9'sd158;
	qsin_lut[6658] =  9'sd62;
	icos_lut[6658] =  9'sd149;
	qsin_lut[6659] =  9'sd89;
	icos_lut[6659] =  9'sd134;
	qsin_lut[6660] =  9'sd114;
	icos_lut[6660] =  9'sd114;
	qsin_lut[6661] =  9'sd134;
	icos_lut[6661] =  9'sd89;
	qsin_lut[6662] =  9'sd149;
	icos_lut[6662] =  9'sd62;
	qsin_lut[6663] =  9'sd158;
	icos_lut[6663] =  9'sd31;
	qsin_lut[6664] =  9'sd161;
	icos_lut[6664] =  9'sd0;
	qsin_lut[6665] =  9'sd158;
	icos_lut[6665] = -9'sd31;
	qsin_lut[6666] =  9'sd149;
	icos_lut[6666] = -9'sd62;
	qsin_lut[6667] =  9'sd134;
	icos_lut[6667] = -9'sd89;
	qsin_lut[6668] =  9'sd114;
	icos_lut[6668] = -9'sd114;
	qsin_lut[6669] =  9'sd89;
	icos_lut[6669] = -9'sd134;
	qsin_lut[6670] =  9'sd62;
	icos_lut[6670] = -9'sd149;
	qsin_lut[6671] =  9'sd31;
	icos_lut[6671] = -9'sd158;
	qsin_lut[6672] =  9'sd0;
	icos_lut[6672] = -9'sd161;
	qsin_lut[6673] = -9'sd31;
	icos_lut[6673] = -9'sd158;
	qsin_lut[6674] = -9'sd62;
	icos_lut[6674] = -9'sd149;
	qsin_lut[6675] = -9'sd89;
	icos_lut[6675] = -9'sd134;
	qsin_lut[6676] = -9'sd114;
	icos_lut[6676] = -9'sd114;
	qsin_lut[6677] = -9'sd134;
	icos_lut[6677] = -9'sd89;
	qsin_lut[6678] = -9'sd149;
	icos_lut[6678] = -9'sd62;
	qsin_lut[6679] = -9'sd158;
	icos_lut[6679] = -9'sd31;
	qsin_lut[6680] = -9'sd161;
	icos_lut[6680] = -9'sd0;
	qsin_lut[6681] = -9'sd158;
	icos_lut[6681] =  9'sd31;
	qsin_lut[6682] = -9'sd149;
	icos_lut[6682] =  9'sd62;
	qsin_lut[6683] = -9'sd134;
	icos_lut[6683] =  9'sd89;
	qsin_lut[6684] = -9'sd114;
	icos_lut[6684] =  9'sd114;
	qsin_lut[6685] = -9'sd89;
	icos_lut[6685] =  9'sd134;
	qsin_lut[6686] = -9'sd62;
	icos_lut[6686] =  9'sd149;
	qsin_lut[6687] = -9'sd31;
	icos_lut[6687] =  9'sd158;
	qsin_lut[6688] =  9'sd0;
	icos_lut[6688] =  9'sd163;
	qsin_lut[6689] =  9'sd32;
	icos_lut[6689] =  9'sd160;
	qsin_lut[6690] =  9'sd62;
	icos_lut[6690] =  9'sd151;
	qsin_lut[6691] =  9'sd91;
	icos_lut[6691] =  9'sd136;
	qsin_lut[6692] =  9'sd115;
	icos_lut[6692] =  9'sd115;
	qsin_lut[6693] =  9'sd136;
	icos_lut[6693] =  9'sd91;
	qsin_lut[6694] =  9'sd151;
	icos_lut[6694] =  9'sd62;
	qsin_lut[6695] =  9'sd160;
	icos_lut[6695] =  9'sd32;
	qsin_lut[6696] =  9'sd163;
	icos_lut[6696] =  9'sd0;
	qsin_lut[6697] =  9'sd160;
	icos_lut[6697] = -9'sd32;
	qsin_lut[6698] =  9'sd151;
	icos_lut[6698] = -9'sd62;
	qsin_lut[6699] =  9'sd136;
	icos_lut[6699] = -9'sd91;
	qsin_lut[6700] =  9'sd115;
	icos_lut[6700] = -9'sd115;
	qsin_lut[6701] =  9'sd91;
	icos_lut[6701] = -9'sd136;
	qsin_lut[6702] =  9'sd62;
	icos_lut[6702] = -9'sd151;
	qsin_lut[6703] =  9'sd32;
	icos_lut[6703] = -9'sd160;
	qsin_lut[6704] =  9'sd0;
	icos_lut[6704] = -9'sd163;
	qsin_lut[6705] = -9'sd32;
	icos_lut[6705] = -9'sd160;
	qsin_lut[6706] = -9'sd62;
	icos_lut[6706] = -9'sd151;
	qsin_lut[6707] = -9'sd91;
	icos_lut[6707] = -9'sd136;
	qsin_lut[6708] = -9'sd115;
	icos_lut[6708] = -9'sd115;
	qsin_lut[6709] = -9'sd136;
	icos_lut[6709] = -9'sd91;
	qsin_lut[6710] = -9'sd151;
	icos_lut[6710] = -9'sd62;
	qsin_lut[6711] = -9'sd160;
	icos_lut[6711] = -9'sd32;
	qsin_lut[6712] = -9'sd163;
	icos_lut[6712] = -9'sd0;
	qsin_lut[6713] = -9'sd160;
	icos_lut[6713] =  9'sd32;
	qsin_lut[6714] = -9'sd151;
	icos_lut[6714] =  9'sd62;
	qsin_lut[6715] = -9'sd136;
	icos_lut[6715] =  9'sd91;
	qsin_lut[6716] = -9'sd115;
	icos_lut[6716] =  9'sd115;
	qsin_lut[6717] = -9'sd91;
	icos_lut[6717] =  9'sd136;
	qsin_lut[6718] = -9'sd62;
	icos_lut[6718] =  9'sd151;
	qsin_lut[6719] = -9'sd32;
	icos_lut[6719] =  9'sd160;
	qsin_lut[6720] =  9'sd0;
	icos_lut[6720] =  9'sd165;
	qsin_lut[6721] =  9'sd32;
	icos_lut[6721] =  9'sd162;
	qsin_lut[6722] =  9'sd63;
	icos_lut[6722] =  9'sd152;
	qsin_lut[6723] =  9'sd92;
	icos_lut[6723] =  9'sd137;
	qsin_lut[6724] =  9'sd117;
	icos_lut[6724] =  9'sd117;
	qsin_lut[6725] =  9'sd137;
	icos_lut[6725] =  9'sd92;
	qsin_lut[6726] =  9'sd152;
	icos_lut[6726] =  9'sd63;
	qsin_lut[6727] =  9'sd162;
	icos_lut[6727] =  9'sd32;
	qsin_lut[6728] =  9'sd165;
	icos_lut[6728] =  9'sd0;
	qsin_lut[6729] =  9'sd162;
	icos_lut[6729] = -9'sd32;
	qsin_lut[6730] =  9'sd152;
	icos_lut[6730] = -9'sd63;
	qsin_lut[6731] =  9'sd137;
	icos_lut[6731] = -9'sd92;
	qsin_lut[6732] =  9'sd117;
	icos_lut[6732] = -9'sd117;
	qsin_lut[6733] =  9'sd92;
	icos_lut[6733] = -9'sd137;
	qsin_lut[6734] =  9'sd63;
	icos_lut[6734] = -9'sd152;
	qsin_lut[6735] =  9'sd32;
	icos_lut[6735] = -9'sd162;
	qsin_lut[6736] =  9'sd0;
	icos_lut[6736] = -9'sd165;
	qsin_lut[6737] = -9'sd32;
	icos_lut[6737] = -9'sd162;
	qsin_lut[6738] = -9'sd63;
	icos_lut[6738] = -9'sd152;
	qsin_lut[6739] = -9'sd92;
	icos_lut[6739] = -9'sd137;
	qsin_lut[6740] = -9'sd117;
	icos_lut[6740] = -9'sd117;
	qsin_lut[6741] = -9'sd137;
	icos_lut[6741] = -9'sd92;
	qsin_lut[6742] = -9'sd152;
	icos_lut[6742] = -9'sd63;
	qsin_lut[6743] = -9'sd162;
	icos_lut[6743] = -9'sd32;
	qsin_lut[6744] = -9'sd165;
	icos_lut[6744] = -9'sd0;
	qsin_lut[6745] = -9'sd162;
	icos_lut[6745] =  9'sd32;
	qsin_lut[6746] = -9'sd152;
	icos_lut[6746] =  9'sd63;
	qsin_lut[6747] = -9'sd137;
	icos_lut[6747] =  9'sd92;
	qsin_lut[6748] = -9'sd117;
	icos_lut[6748] =  9'sd117;
	qsin_lut[6749] = -9'sd92;
	icos_lut[6749] =  9'sd137;
	qsin_lut[6750] = -9'sd63;
	icos_lut[6750] =  9'sd152;
	qsin_lut[6751] = -9'sd32;
	icos_lut[6751] =  9'sd162;
	qsin_lut[6752] =  9'sd0;
	icos_lut[6752] =  9'sd167;
	qsin_lut[6753] =  9'sd33;
	icos_lut[6753] =  9'sd164;
	qsin_lut[6754] =  9'sd64;
	icos_lut[6754] =  9'sd154;
	qsin_lut[6755] =  9'sd93;
	icos_lut[6755] =  9'sd139;
	qsin_lut[6756] =  9'sd118;
	icos_lut[6756] =  9'sd118;
	qsin_lut[6757] =  9'sd139;
	icos_lut[6757] =  9'sd93;
	qsin_lut[6758] =  9'sd154;
	icos_lut[6758] =  9'sd64;
	qsin_lut[6759] =  9'sd164;
	icos_lut[6759] =  9'sd33;
	qsin_lut[6760] =  9'sd167;
	icos_lut[6760] =  9'sd0;
	qsin_lut[6761] =  9'sd164;
	icos_lut[6761] = -9'sd33;
	qsin_lut[6762] =  9'sd154;
	icos_lut[6762] = -9'sd64;
	qsin_lut[6763] =  9'sd139;
	icos_lut[6763] = -9'sd93;
	qsin_lut[6764] =  9'sd118;
	icos_lut[6764] = -9'sd118;
	qsin_lut[6765] =  9'sd93;
	icos_lut[6765] = -9'sd139;
	qsin_lut[6766] =  9'sd64;
	icos_lut[6766] = -9'sd154;
	qsin_lut[6767] =  9'sd33;
	icos_lut[6767] = -9'sd164;
	qsin_lut[6768] =  9'sd0;
	icos_lut[6768] = -9'sd167;
	qsin_lut[6769] = -9'sd33;
	icos_lut[6769] = -9'sd164;
	qsin_lut[6770] = -9'sd64;
	icos_lut[6770] = -9'sd154;
	qsin_lut[6771] = -9'sd93;
	icos_lut[6771] = -9'sd139;
	qsin_lut[6772] = -9'sd118;
	icos_lut[6772] = -9'sd118;
	qsin_lut[6773] = -9'sd139;
	icos_lut[6773] = -9'sd93;
	qsin_lut[6774] = -9'sd154;
	icos_lut[6774] = -9'sd64;
	qsin_lut[6775] = -9'sd164;
	icos_lut[6775] = -9'sd33;
	qsin_lut[6776] = -9'sd167;
	icos_lut[6776] = -9'sd0;
	qsin_lut[6777] = -9'sd164;
	icos_lut[6777] =  9'sd33;
	qsin_lut[6778] = -9'sd154;
	icos_lut[6778] =  9'sd64;
	qsin_lut[6779] = -9'sd139;
	icos_lut[6779] =  9'sd93;
	qsin_lut[6780] = -9'sd118;
	icos_lut[6780] =  9'sd118;
	qsin_lut[6781] = -9'sd93;
	icos_lut[6781] =  9'sd139;
	qsin_lut[6782] = -9'sd64;
	icos_lut[6782] =  9'sd154;
	qsin_lut[6783] = -9'sd33;
	icos_lut[6783] =  9'sd164;
	qsin_lut[6784] =  9'sd0;
	icos_lut[6784] =  9'sd169;
	qsin_lut[6785] =  9'sd33;
	icos_lut[6785] =  9'sd166;
	qsin_lut[6786] =  9'sd65;
	icos_lut[6786] =  9'sd156;
	qsin_lut[6787] =  9'sd94;
	icos_lut[6787] =  9'sd141;
	qsin_lut[6788] =  9'sd120;
	icos_lut[6788] =  9'sd120;
	qsin_lut[6789] =  9'sd141;
	icos_lut[6789] =  9'sd94;
	qsin_lut[6790] =  9'sd156;
	icos_lut[6790] =  9'sd65;
	qsin_lut[6791] =  9'sd166;
	icos_lut[6791] =  9'sd33;
	qsin_lut[6792] =  9'sd169;
	icos_lut[6792] =  9'sd0;
	qsin_lut[6793] =  9'sd166;
	icos_lut[6793] = -9'sd33;
	qsin_lut[6794] =  9'sd156;
	icos_lut[6794] = -9'sd65;
	qsin_lut[6795] =  9'sd141;
	icos_lut[6795] = -9'sd94;
	qsin_lut[6796] =  9'sd120;
	icos_lut[6796] = -9'sd120;
	qsin_lut[6797] =  9'sd94;
	icos_lut[6797] = -9'sd141;
	qsin_lut[6798] =  9'sd65;
	icos_lut[6798] = -9'sd156;
	qsin_lut[6799] =  9'sd33;
	icos_lut[6799] = -9'sd166;
	qsin_lut[6800] =  9'sd0;
	icos_lut[6800] = -9'sd169;
	qsin_lut[6801] = -9'sd33;
	icos_lut[6801] = -9'sd166;
	qsin_lut[6802] = -9'sd65;
	icos_lut[6802] = -9'sd156;
	qsin_lut[6803] = -9'sd94;
	icos_lut[6803] = -9'sd141;
	qsin_lut[6804] = -9'sd120;
	icos_lut[6804] = -9'sd120;
	qsin_lut[6805] = -9'sd141;
	icos_lut[6805] = -9'sd94;
	qsin_lut[6806] = -9'sd156;
	icos_lut[6806] = -9'sd65;
	qsin_lut[6807] = -9'sd166;
	icos_lut[6807] = -9'sd33;
	qsin_lut[6808] = -9'sd169;
	icos_lut[6808] = -9'sd0;
	qsin_lut[6809] = -9'sd166;
	icos_lut[6809] =  9'sd33;
	qsin_lut[6810] = -9'sd156;
	icos_lut[6810] =  9'sd65;
	qsin_lut[6811] = -9'sd141;
	icos_lut[6811] =  9'sd94;
	qsin_lut[6812] = -9'sd120;
	icos_lut[6812] =  9'sd120;
	qsin_lut[6813] = -9'sd94;
	icos_lut[6813] =  9'sd141;
	qsin_lut[6814] = -9'sd65;
	icos_lut[6814] =  9'sd156;
	qsin_lut[6815] = -9'sd33;
	icos_lut[6815] =  9'sd166;
	qsin_lut[6816] =  9'sd0;
	icos_lut[6816] =  9'sd171;
	qsin_lut[6817] =  9'sd33;
	icos_lut[6817] =  9'sd168;
	qsin_lut[6818] =  9'sd65;
	icos_lut[6818] =  9'sd158;
	qsin_lut[6819] =  9'sd95;
	icos_lut[6819] =  9'sd142;
	qsin_lut[6820] =  9'sd121;
	icos_lut[6820] =  9'sd121;
	qsin_lut[6821] =  9'sd142;
	icos_lut[6821] =  9'sd95;
	qsin_lut[6822] =  9'sd158;
	icos_lut[6822] =  9'sd65;
	qsin_lut[6823] =  9'sd168;
	icos_lut[6823] =  9'sd33;
	qsin_lut[6824] =  9'sd171;
	icos_lut[6824] =  9'sd0;
	qsin_lut[6825] =  9'sd168;
	icos_lut[6825] = -9'sd33;
	qsin_lut[6826] =  9'sd158;
	icos_lut[6826] = -9'sd65;
	qsin_lut[6827] =  9'sd142;
	icos_lut[6827] = -9'sd95;
	qsin_lut[6828] =  9'sd121;
	icos_lut[6828] = -9'sd121;
	qsin_lut[6829] =  9'sd95;
	icos_lut[6829] = -9'sd142;
	qsin_lut[6830] =  9'sd65;
	icos_lut[6830] = -9'sd158;
	qsin_lut[6831] =  9'sd33;
	icos_lut[6831] = -9'sd168;
	qsin_lut[6832] =  9'sd0;
	icos_lut[6832] = -9'sd171;
	qsin_lut[6833] = -9'sd33;
	icos_lut[6833] = -9'sd168;
	qsin_lut[6834] = -9'sd65;
	icos_lut[6834] = -9'sd158;
	qsin_lut[6835] = -9'sd95;
	icos_lut[6835] = -9'sd142;
	qsin_lut[6836] = -9'sd121;
	icos_lut[6836] = -9'sd121;
	qsin_lut[6837] = -9'sd142;
	icos_lut[6837] = -9'sd95;
	qsin_lut[6838] = -9'sd158;
	icos_lut[6838] = -9'sd65;
	qsin_lut[6839] = -9'sd168;
	icos_lut[6839] = -9'sd33;
	qsin_lut[6840] = -9'sd171;
	icos_lut[6840] = -9'sd0;
	qsin_lut[6841] = -9'sd168;
	icos_lut[6841] =  9'sd33;
	qsin_lut[6842] = -9'sd158;
	icos_lut[6842] =  9'sd65;
	qsin_lut[6843] = -9'sd142;
	icos_lut[6843] =  9'sd95;
	qsin_lut[6844] = -9'sd121;
	icos_lut[6844] =  9'sd121;
	qsin_lut[6845] = -9'sd95;
	icos_lut[6845] =  9'sd142;
	qsin_lut[6846] = -9'sd65;
	icos_lut[6846] =  9'sd158;
	qsin_lut[6847] = -9'sd33;
	icos_lut[6847] =  9'sd168;
	qsin_lut[6848] =  9'sd0;
	icos_lut[6848] =  9'sd173;
	qsin_lut[6849] =  9'sd34;
	icos_lut[6849] =  9'sd170;
	qsin_lut[6850] =  9'sd66;
	icos_lut[6850] =  9'sd160;
	qsin_lut[6851] =  9'sd96;
	icos_lut[6851] =  9'sd144;
	qsin_lut[6852] =  9'sd122;
	icos_lut[6852] =  9'sd122;
	qsin_lut[6853] =  9'sd144;
	icos_lut[6853] =  9'sd96;
	qsin_lut[6854] =  9'sd160;
	icos_lut[6854] =  9'sd66;
	qsin_lut[6855] =  9'sd170;
	icos_lut[6855] =  9'sd34;
	qsin_lut[6856] =  9'sd173;
	icos_lut[6856] =  9'sd0;
	qsin_lut[6857] =  9'sd170;
	icos_lut[6857] = -9'sd34;
	qsin_lut[6858] =  9'sd160;
	icos_lut[6858] = -9'sd66;
	qsin_lut[6859] =  9'sd144;
	icos_lut[6859] = -9'sd96;
	qsin_lut[6860] =  9'sd122;
	icos_lut[6860] = -9'sd122;
	qsin_lut[6861] =  9'sd96;
	icos_lut[6861] = -9'sd144;
	qsin_lut[6862] =  9'sd66;
	icos_lut[6862] = -9'sd160;
	qsin_lut[6863] =  9'sd34;
	icos_lut[6863] = -9'sd170;
	qsin_lut[6864] =  9'sd0;
	icos_lut[6864] = -9'sd173;
	qsin_lut[6865] = -9'sd34;
	icos_lut[6865] = -9'sd170;
	qsin_lut[6866] = -9'sd66;
	icos_lut[6866] = -9'sd160;
	qsin_lut[6867] = -9'sd96;
	icos_lut[6867] = -9'sd144;
	qsin_lut[6868] = -9'sd122;
	icos_lut[6868] = -9'sd122;
	qsin_lut[6869] = -9'sd144;
	icos_lut[6869] = -9'sd96;
	qsin_lut[6870] = -9'sd160;
	icos_lut[6870] = -9'sd66;
	qsin_lut[6871] = -9'sd170;
	icos_lut[6871] = -9'sd34;
	qsin_lut[6872] = -9'sd173;
	icos_lut[6872] = -9'sd0;
	qsin_lut[6873] = -9'sd170;
	icos_lut[6873] =  9'sd34;
	qsin_lut[6874] = -9'sd160;
	icos_lut[6874] =  9'sd66;
	qsin_lut[6875] = -9'sd144;
	icos_lut[6875] =  9'sd96;
	qsin_lut[6876] = -9'sd122;
	icos_lut[6876] =  9'sd122;
	qsin_lut[6877] = -9'sd96;
	icos_lut[6877] =  9'sd144;
	qsin_lut[6878] = -9'sd66;
	icos_lut[6878] =  9'sd160;
	qsin_lut[6879] = -9'sd34;
	icos_lut[6879] =  9'sd170;
	qsin_lut[6880] =  9'sd0;
	icos_lut[6880] =  9'sd175;
	qsin_lut[6881] =  9'sd34;
	icos_lut[6881] =  9'sd172;
	qsin_lut[6882] =  9'sd67;
	icos_lut[6882] =  9'sd162;
	qsin_lut[6883] =  9'sd97;
	icos_lut[6883] =  9'sd146;
	qsin_lut[6884] =  9'sd124;
	icos_lut[6884] =  9'sd124;
	qsin_lut[6885] =  9'sd146;
	icos_lut[6885] =  9'sd97;
	qsin_lut[6886] =  9'sd162;
	icos_lut[6886] =  9'sd67;
	qsin_lut[6887] =  9'sd172;
	icos_lut[6887] =  9'sd34;
	qsin_lut[6888] =  9'sd175;
	icos_lut[6888] =  9'sd0;
	qsin_lut[6889] =  9'sd172;
	icos_lut[6889] = -9'sd34;
	qsin_lut[6890] =  9'sd162;
	icos_lut[6890] = -9'sd67;
	qsin_lut[6891] =  9'sd146;
	icos_lut[6891] = -9'sd97;
	qsin_lut[6892] =  9'sd124;
	icos_lut[6892] = -9'sd124;
	qsin_lut[6893] =  9'sd97;
	icos_lut[6893] = -9'sd146;
	qsin_lut[6894] =  9'sd67;
	icos_lut[6894] = -9'sd162;
	qsin_lut[6895] =  9'sd34;
	icos_lut[6895] = -9'sd172;
	qsin_lut[6896] =  9'sd0;
	icos_lut[6896] = -9'sd175;
	qsin_lut[6897] = -9'sd34;
	icos_lut[6897] = -9'sd172;
	qsin_lut[6898] = -9'sd67;
	icos_lut[6898] = -9'sd162;
	qsin_lut[6899] = -9'sd97;
	icos_lut[6899] = -9'sd146;
	qsin_lut[6900] = -9'sd124;
	icos_lut[6900] = -9'sd124;
	qsin_lut[6901] = -9'sd146;
	icos_lut[6901] = -9'sd97;
	qsin_lut[6902] = -9'sd162;
	icos_lut[6902] = -9'sd67;
	qsin_lut[6903] = -9'sd172;
	icos_lut[6903] = -9'sd34;
	qsin_lut[6904] = -9'sd175;
	icos_lut[6904] = -9'sd0;
	qsin_lut[6905] = -9'sd172;
	icos_lut[6905] =  9'sd34;
	qsin_lut[6906] = -9'sd162;
	icos_lut[6906] =  9'sd67;
	qsin_lut[6907] = -9'sd146;
	icos_lut[6907] =  9'sd97;
	qsin_lut[6908] = -9'sd124;
	icos_lut[6908] =  9'sd124;
	qsin_lut[6909] = -9'sd97;
	icos_lut[6909] =  9'sd146;
	qsin_lut[6910] = -9'sd67;
	icos_lut[6910] =  9'sd162;
	qsin_lut[6911] = -9'sd34;
	icos_lut[6911] =  9'sd172;
	qsin_lut[6912] =  9'sd0;
	icos_lut[6912] =  9'sd177;
	qsin_lut[6913] =  9'sd35;
	icos_lut[6913] =  9'sd174;
	qsin_lut[6914] =  9'sd68;
	icos_lut[6914] =  9'sd164;
	qsin_lut[6915] =  9'sd98;
	icos_lut[6915] =  9'sd147;
	qsin_lut[6916] =  9'sd125;
	icos_lut[6916] =  9'sd125;
	qsin_lut[6917] =  9'sd147;
	icos_lut[6917] =  9'sd98;
	qsin_lut[6918] =  9'sd164;
	icos_lut[6918] =  9'sd68;
	qsin_lut[6919] =  9'sd174;
	icos_lut[6919] =  9'sd35;
	qsin_lut[6920] =  9'sd177;
	icos_lut[6920] =  9'sd0;
	qsin_lut[6921] =  9'sd174;
	icos_lut[6921] = -9'sd35;
	qsin_lut[6922] =  9'sd164;
	icos_lut[6922] = -9'sd68;
	qsin_lut[6923] =  9'sd147;
	icos_lut[6923] = -9'sd98;
	qsin_lut[6924] =  9'sd125;
	icos_lut[6924] = -9'sd125;
	qsin_lut[6925] =  9'sd98;
	icos_lut[6925] = -9'sd147;
	qsin_lut[6926] =  9'sd68;
	icos_lut[6926] = -9'sd164;
	qsin_lut[6927] =  9'sd35;
	icos_lut[6927] = -9'sd174;
	qsin_lut[6928] =  9'sd0;
	icos_lut[6928] = -9'sd177;
	qsin_lut[6929] = -9'sd35;
	icos_lut[6929] = -9'sd174;
	qsin_lut[6930] = -9'sd68;
	icos_lut[6930] = -9'sd164;
	qsin_lut[6931] = -9'sd98;
	icos_lut[6931] = -9'sd147;
	qsin_lut[6932] = -9'sd125;
	icos_lut[6932] = -9'sd125;
	qsin_lut[6933] = -9'sd147;
	icos_lut[6933] = -9'sd98;
	qsin_lut[6934] = -9'sd164;
	icos_lut[6934] = -9'sd68;
	qsin_lut[6935] = -9'sd174;
	icos_lut[6935] = -9'sd35;
	qsin_lut[6936] = -9'sd177;
	icos_lut[6936] = -9'sd0;
	qsin_lut[6937] = -9'sd174;
	icos_lut[6937] =  9'sd35;
	qsin_lut[6938] = -9'sd164;
	icos_lut[6938] =  9'sd68;
	qsin_lut[6939] = -9'sd147;
	icos_lut[6939] =  9'sd98;
	qsin_lut[6940] = -9'sd125;
	icos_lut[6940] =  9'sd125;
	qsin_lut[6941] = -9'sd98;
	icos_lut[6941] =  9'sd147;
	qsin_lut[6942] = -9'sd68;
	icos_lut[6942] =  9'sd164;
	qsin_lut[6943] = -9'sd35;
	icos_lut[6943] =  9'sd174;
	qsin_lut[6944] =  9'sd0;
	icos_lut[6944] =  9'sd179;
	qsin_lut[6945] =  9'sd35;
	icos_lut[6945] =  9'sd176;
	qsin_lut[6946] =  9'sd69;
	icos_lut[6946] =  9'sd165;
	qsin_lut[6947] =  9'sd99;
	icos_lut[6947] =  9'sd149;
	qsin_lut[6948] =  9'sd127;
	icos_lut[6948] =  9'sd127;
	qsin_lut[6949] =  9'sd149;
	icos_lut[6949] =  9'sd99;
	qsin_lut[6950] =  9'sd165;
	icos_lut[6950] =  9'sd69;
	qsin_lut[6951] =  9'sd176;
	icos_lut[6951] =  9'sd35;
	qsin_lut[6952] =  9'sd179;
	icos_lut[6952] =  9'sd0;
	qsin_lut[6953] =  9'sd176;
	icos_lut[6953] = -9'sd35;
	qsin_lut[6954] =  9'sd165;
	icos_lut[6954] = -9'sd69;
	qsin_lut[6955] =  9'sd149;
	icos_lut[6955] = -9'sd99;
	qsin_lut[6956] =  9'sd127;
	icos_lut[6956] = -9'sd127;
	qsin_lut[6957] =  9'sd99;
	icos_lut[6957] = -9'sd149;
	qsin_lut[6958] =  9'sd69;
	icos_lut[6958] = -9'sd165;
	qsin_lut[6959] =  9'sd35;
	icos_lut[6959] = -9'sd176;
	qsin_lut[6960] =  9'sd0;
	icos_lut[6960] = -9'sd179;
	qsin_lut[6961] = -9'sd35;
	icos_lut[6961] = -9'sd176;
	qsin_lut[6962] = -9'sd69;
	icos_lut[6962] = -9'sd165;
	qsin_lut[6963] = -9'sd99;
	icos_lut[6963] = -9'sd149;
	qsin_lut[6964] = -9'sd127;
	icos_lut[6964] = -9'sd127;
	qsin_lut[6965] = -9'sd149;
	icos_lut[6965] = -9'sd99;
	qsin_lut[6966] = -9'sd165;
	icos_lut[6966] = -9'sd69;
	qsin_lut[6967] = -9'sd176;
	icos_lut[6967] = -9'sd35;
	qsin_lut[6968] = -9'sd179;
	icos_lut[6968] = -9'sd0;
	qsin_lut[6969] = -9'sd176;
	icos_lut[6969] =  9'sd35;
	qsin_lut[6970] = -9'sd165;
	icos_lut[6970] =  9'sd69;
	qsin_lut[6971] = -9'sd149;
	icos_lut[6971] =  9'sd99;
	qsin_lut[6972] = -9'sd127;
	icos_lut[6972] =  9'sd127;
	qsin_lut[6973] = -9'sd99;
	icos_lut[6973] =  9'sd149;
	qsin_lut[6974] = -9'sd69;
	icos_lut[6974] =  9'sd165;
	qsin_lut[6975] = -9'sd35;
	icos_lut[6975] =  9'sd176;
	qsin_lut[6976] =  9'sd0;
	icos_lut[6976] =  9'sd181;
	qsin_lut[6977] =  9'sd35;
	icos_lut[6977] =  9'sd178;
	qsin_lut[6978] =  9'sd69;
	icos_lut[6978] =  9'sd167;
	qsin_lut[6979] =  9'sd101;
	icos_lut[6979] =  9'sd150;
	qsin_lut[6980] =  9'sd128;
	icos_lut[6980] =  9'sd128;
	qsin_lut[6981] =  9'sd150;
	icos_lut[6981] =  9'sd101;
	qsin_lut[6982] =  9'sd167;
	icos_lut[6982] =  9'sd69;
	qsin_lut[6983] =  9'sd178;
	icos_lut[6983] =  9'sd35;
	qsin_lut[6984] =  9'sd181;
	icos_lut[6984] =  9'sd0;
	qsin_lut[6985] =  9'sd178;
	icos_lut[6985] = -9'sd35;
	qsin_lut[6986] =  9'sd167;
	icos_lut[6986] = -9'sd69;
	qsin_lut[6987] =  9'sd150;
	icos_lut[6987] = -9'sd101;
	qsin_lut[6988] =  9'sd128;
	icos_lut[6988] = -9'sd128;
	qsin_lut[6989] =  9'sd101;
	icos_lut[6989] = -9'sd150;
	qsin_lut[6990] =  9'sd69;
	icos_lut[6990] = -9'sd167;
	qsin_lut[6991] =  9'sd35;
	icos_lut[6991] = -9'sd178;
	qsin_lut[6992] =  9'sd0;
	icos_lut[6992] = -9'sd181;
	qsin_lut[6993] = -9'sd35;
	icos_lut[6993] = -9'sd178;
	qsin_lut[6994] = -9'sd69;
	icos_lut[6994] = -9'sd167;
	qsin_lut[6995] = -9'sd101;
	icos_lut[6995] = -9'sd150;
	qsin_lut[6996] = -9'sd128;
	icos_lut[6996] = -9'sd128;
	qsin_lut[6997] = -9'sd150;
	icos_lut[6997] = -9'sd101;
	qsin_lut[6998] = -9'sd167;
	icos_lut[6998] = -9'sd69;
	qsin_lut[6999] = -9'sd178;
	icos_lut[6999] = -9'sd35;
	qsin_lut[7000] = -9'sd181;
	icos_lut[7000] = -9'sd0;
	qsin_lut[7001] = -9'sd178;
	icos_lut[7001] =  9'sd35;
	qsin_lut[7002] = -9'sd167;
	icos_lut[7002] =  9'sd69;
	qsin_lut[7003] = -9'sd150;
	icos_lut[7003] =  9'sd101;
	qsin_lut[7004] = -9'sd128;
	icos_lut[7004] =  9'sd128;
	qsin_lut[7005] = -9'sd101;
	icos_lut[7005] =  9'sd150;
	qsin_lut[7006] = -9'sd69;
	icos_lut[7006] =  9'sd167;
	qsin_lut[7007] = -9'sd35;
	icos_lut[7007] =  9'sd178;
	qsin_lut[7008] =  9'sd0;
	icos_lut[7008] =  9'sd183;
	qsin_lut[7009] =  9'sd36;
	icos_lut[7009] =  9'sd179;
	qsin_lut[7010] =  9'sd70;
	icos_lut[7010] =  9'sd169;
	qsin_lut[7011] =  9'sd102;
	icos_lut[7011] =  9'sd152;
	qsin_lut[7012] =  9'sd129;
	icos_lut[7012] =  9'sd129;
	qsin_lut[7013] =  9'sd152;
	icos_lut[7013] =  9'sd102;
	qsin_lut[7014] =  9'sd169;
	icos_lut[7014] =  9'sd70;
	qsin_lut[7015] =  9'sd179;
	icos_lut[7015] =  9'sd36;
	qsin_lut[7016] =  9'sd183;
	icos_lut[7016] =  9'sd0;
	qsin_lut[7017] =  9'sd179;
	icos_lut[7017] = -9'sd36;
	qsin_lut[7018] =  9'sd169;
	icos_lut[7018] = -9'sd70;
	qsin_lut[7019] =  9'sd152;
	icos_lut[7019] = -9'sd102;
	qsin_lut[7020] =  9'sd129;
	icos_lut[7020] = -9'sd129;
	qsin_lut[7021] =  9'sd102;
	icos_lut[7021] = -9'sd152;
	qsin_lut[7022] =  9'sd70;
	icos_lut[7022] = -9'sd169;
	qsin_lut[7023] =  9'sd36;
	icos_lut[7023] = -9'sd179;
	qsin_lut[7024] =  9'sd0;
	icos_lut[7024] = -9'sd183;
	qsin_lut[7025] = -9'sd36;
	icos_lut[7025] = -9'sd179;
	qsin_lut[7026] = -9'sd70;
	icos_lut[7026] = -9'sd169;
	qsin_lut[7027] = -9'sd102;
	icos_lut[7027] = -9'sd152;
	qsin_lut[7028] = -9'sd129;
	icos_lut[7028] = -9'sd129;
	qsin_lut[7029] = -9'sd152;
	icos_lut[7029] = -9'sd102;
	qsin_lut[7030] = -9'sd169;
	icos_lut[7030] = -9'sd70;
	qsin_lut[7031] = -9'sd179;
	icos_lut[7031] = -9'sd36;
	qsin_lut[7032] = -9'sd183;
	icos_lut[7032] = -9'sd0;
	qsin_lut[7033] = -9'sd179;
	icos_lut[7033] =  9'sd36;
	qsin_lut[7034] = -9'sd169;
	icos_lut[7034] =  9'sd70;
	qsin_lut[7035] = -9'sd152;
	icos_lut[7035] =  9'sd102;
	qsin_lut[7036] = -9'sd129;
	icos_lut[7036] =  9'sd129;
	qsin_lut[7037] = -9'sd102;
	icos_lut[7037] =  9'sd152;
	qsin_lut[7038] = -9'sd70;
	icos_lut[7038] =  9'sd169;
	qsin_lut[7039] = -9'sd36;
	icos_lut[7039] =  9'sd179;
	qsin_lut[7040] =  9'sd0;
	icos_lut[7040] =  9'sd185;
	qsin_lut[7041] =  9'sd36;
	icos_lut[7041] =  9'sd181;
	qsin_lut[7042] =  9'sd71;
	icos_lut[7042] =  9'sd171;
	qsin_lut[7043] =  9'sd103;
	icos_lut[7043] =  9'sd154;
	qsin_lut[7044] =  9'sd131;
	icos_lut[7044] =  9'sd131;
	qsin_lut[7045] =  9'sd154;
	icos_lut[7045] =  9'sd103;
	qsin_lut[7046] =  9'sd171;
	icos_lut[7046] =  9'sd71;
	qsin_lut[7047] =  9'sd181;
	icos_lut[7047] =  9'sd36;
	qsin_lut[7048] =  9'sd185;
	icos_lut[7048] =  9'sd0;
	qsin_lut[7049] =  9'sd181;
	icos_lut[7049] = -9'sd36;
	qsin_lut[7050] =  9'sd171;
	icos_lut[7050] = -9'sd71;
	qsin_lut[7051] =  9'sd154;
	icos_lut[7051] = -9'sd103;
	qsin_lut[7052] =  9'sd131;
	icos_lut[7052] = -9'sd131;
	qsin_lut[7053] =  9'sd103;
	icos_lut[7053] = -9'sd154;
	qsin_lut[7054] =  9'sd71;
	icos_lut[7054] = -9'sd171;
	qsin_lut[7055] =  9'sd36;
	icos_lut[7055] = -9'sd181;
	qsin_lut[7056] =  9'sd0;
	icos_lut[7056] = -9'sd185;
	qsin_lut[7057] = -9'sd36;
	icos_lut[7057] = -9'sd181;
	qsin_lut[7058] = -9'sd71;
	icos_lut[7058] = -9'sd171;
	qsin_lut[7059] = -9'sd103;
	icos_lut[7059] = -9'sd154;
	qsin_lut[7060] = -9'sd131;
	icos_lut[7060] = -9'sd131;
	qsin_lut[7061] = -9'sd154;
	icos_lut[7061] = -9'sd103;
	qsin_lut[7062] = -9'sd171;
	icos_lut[7062] = -9'sd71;
	qsin_lut[7063] = -9'sd181;
	icos_lut[7063] = -9'sd36;
	qsin_lut[7064] = -9'sd185;
	icos_lut[7064] = -9'sd0;
	qsin_lut[7065] = -9'sd181;
	icos_lut[7065] =  9'sd36;
	qsin_lut[7066] = -9'sd171;
	icos_lut[7066] =  9'sd71;
	qsin_lut[7067] = -9'sd154;
	icos_lut[7067] =  9'sd103;
	qsin_lut[7068] = -9'sd131;
	icos_lut[7068] =  9'sd131;
	qsin_lut[7069] = -9'sd103;
	icos_lut[7069] =  9'sd154;
	qsin_lut[7070] = -9'sd71;
	icos_lut[7070] =  9'sd171;
	qsin_lut[7071] = -9'sd36;
	icos_lut[7071] =  9'sd181;
	qsin_lut[7072] =  9'sd0;
	icos_lut[7072] =  9'sd187;
	qsin_lut[7073] =  9'sd36;
	icos_lut[7073] =  9'sd183;
	qsin_lut[7074] =  9'sd72;
	icos_lut[7074] =  9'sd173;
	qsin_lut[7075] =  9'sd104;
	icos_lut[7075] =  9'sd155;
	qsin_lut[7076] =  9'sd132;
	icos_lut[7076] =  9'sd132;
	qsin_lut[7077] =  9'sd155;
	icos_lut[7077] =  9'sd104;
	qsin_lut[7078] =  9'sd173;
	icos_lut[7078] =  9'sd72;
	qsin_lut[7079] =  9'sd183;
	icos_lut[7079] =  9'sd36;
	qsin_lut[7080] =  9'sd187;
	icos_lut[7080] =  9'sd0;
	qsin_lut[7081] =  9'sd183;
	icos_lut[7081] = -9'sd36;
	qsin_lut[7082] =  9'sd173;
	icos_lut[7082] = -9'sd72;
	qsin_lut[7083] =  9'sd155;
	icos_lut[7083] = -9'sd104;
	qsin_lut[7084] =  9'sd132;
	icos_lut[7084] = -9'sd132;
	qsin_lut[7085] =  9'sd104;
	icos_lut[7085] = -9'sd155;
	qsin_lut[7086] =  9'sd72;
	icos_lut[7086] = -9'sd173;
	qsin_lut[7087] =  9'sd36;
	icos_lut[7087] = -9'sd183;
	qsin_lut[7088] =  9'sd0;
	icos_lut[7088] = -9'sd187;
	qsin_lut[7089] = -9'sd36;
	icos_lut[7089] = -9'sd183;
	qsin_lut[7090] = -9'sd72;
	icos_lut[7090] = -9'sd173;
	qsin_lut[7091] = -9'sd104;
	icos_lut[7091] = -9'sd155;
	qsin_lut[7092] = -9'sd132;
	icos_lut[7092] = -9'sd132;
	qsin_lut[7093] = -9'sd155;
	icos_lut[7093] = -9'sd104;
	qsin_lut[7094] = -9'sd173;
	icos_lut[7094] = -9'sd72;
	qsin_lut[7095] = -9'sd183;
	icos_lut[7095] = -9'sd36;
	qsin_lut[7096] = -9'sd187;
	icos_lut[7096] = -9'sd0;
	qsin_lut[7097] = -9'sd183;
	icos_lut[7097] =  9'sd36;
	qsin_lut[7098] = -9'sd173;
	icos_lut[7098] =  9'sd72;
	qsin_lut[7099] = -9'sd155;
	icos_lut[7099] =  9'sd104;
	qsin_lut[7100] = -9'sd132;
	icos_lut[7100] =  9'sd132;
	qsin_lut[7101] = -9'sd104;
	icos_lut[7101] =  9'sd155;
	qsin_lut[7102] = -9'sd72;
	icos_lut[7102] =  9'sd173;
	qsin_lut[7103] = -9'sd36;
	icos_lut[7103] =  9'sd183;
	qsin_lut[7104] =  9'sd0;
	icos_lut[7104] =  9'sd189;
	qsin_lut[7105] =  9'sd37;
	icos_lut[7105] =  9'sd185;
	qsin_lut[7106] =  9'sd72;
	icos_lut[7106] =  9'sd175;
	qsin_lut[7107] =  9'sd105;
	icos_lut[7107] =  9'sd157;
	qsin_lut[7108] =  9'sd134;
	icos_lut[7108] =  9'sd134;
	qsin_lut[7109] =  9'sd157;
	icos_lut[7109] =  9'sd105;
	qsin_lut[7110] =  9'sd175;
	icos_lut[7110] =  9'sd72;
	qsin_lut[7111] =  9'sd185;
	icos_lut[7111] =  9'sd37;
	qsin_lut[7112] =  9'sd189;
	icos_lut[7112] =  9'sd0;
	qsin_lut[7113] =  9'sd185;
	icos_lut[7113] = -9'sd37;
	qsin_lut[7114] =  9'sd175;
	icos_lut[7114] = -9'sd72;
	qsin_lut[7115] =  9'sd157;
	icos_lut[7115] = -9'sd105;
	qsin_lut[7116] =  9'sd134;
	icos_lut[7116] = -9'sd134;
	qsin_lut[7117] =  9'sd105;
	icos_lut[7117] = -9'sd157;
	qsin_lut[7118] =  9'sd72;
	icos_lut[7118] = -9'sd175;
	qsin_lut[7119] =  9'sd37;
	icos_lut[7119] = -9'sd185;
	qsin_lut[7120] =  9'sd0;
	icos_lut[7120] = -9'sd189;
	qsin_lut[7121] = -9'sd37;
	icos_lut[7121] = -9'sd185;
	qsin_lut[7122] = -9'sd72;
	icos_lut[7122] = -9'sd175;
	qsin_lut[7123] = -9'sd105;
	icos_lut[7123] = -9'sd157;
	qsin_lut[7124] = -9'sd134;
	icos_lut[7124] = -9'sd134;
	qsin_lut[7125] = -9'sd157;
	icos_lut[7125] = -9'sd105;
	qsin_lut[7126] = -9'sd175;
	icos_lut[7126] = -9'sd72;
	qsin_lut[7127] = -9'sd185;
	icos_lut[7127] = -9'sd37;
	qsin_lut[7128] = -9'sd189;
	icos_lut[7128] = -9'sd0;
	qsin_lut[7129] = -9'sd185;
	icos_lut[7129] =  9'sd37;
	qsin_lut[7130] = -9'sd175;
	icos_lut[7130] =  9'sd72;
	qsin_lut[7131] = -9'sd157;
	icos_lut[7131] =  9'sd105;
	qsin_lut[7132] = -9'sd134;
	icos_lut[7132] =  9'sd134;
	qsin_lut[7133] = -9'sd105;
	icos_lut[7133] =  9'sd157;
	qsin_lut[7134] = -9'sd72;
	icos_lut[7134] =  9'sd175;
	qsin_lut[7135] = -9'sd37;
	icos_lut[7135] =  9'sd185;
	qsin_lut[7136] =  9'sd0;
	icos_lut[7136] =  9'sd191;
	qsin_lut[7137] =  9'sd37;
	icos_lut[7137] =  9'sd187;
	qsin_lut[7138] =  9'sd73;
	icos_lut[7138] =  9'sd176;
	qsin_lut[7139] =  9'sd106;
	icos_lut[7139] =  9'sd159;
	qsin_lut[7140] =  9'sd135;
	icos_lut[7140] =  9'sd135;
	qsin_lut[7141] =  9'sd159;
	icos_lut[7141] =  9'sd106;
	qsin_lut[7142] =  9'sd176;
	icos_lut[7142] =  9'sd73;
	qsin_lut[7143] =  9'sd187;
	icos_lut[7143] =  9'sd37;
	qsin_lut[7144] =  9'sd191;
	icos_lut[7144] =  9'sd0;
	qsin_lut[7145] =  9'sd187;
	icos_lut[7145] = -9'sd37;
	qsin_lut[7146] =  9'sd176;
	icos_lut[7146] = -9'sd73;
	qsin_lut[7147] =  9'sd159;
	icos_lut[7147] = -9'sd106;
	qsin_lut[7148] =  9'sd135;
	icos_lut[7148] = -9'sd135;
	qsin_lut[7149] =  9'sd106;
	icos_lut[7149] = -9'sd159;
	qsin_lut[7150] =  9'sd73;
	icos_lut[7150] = -9'sd176;
	qsin_lut[7151] =  9'sd37;
	icos_lut[7151] = -9'sd187;
	qsin_lut[7152] =  9'sd0;
	icos_lut[7152] = -9'sd191;
	qsin_lut[7153] = -9'sd37;
	icos_lut[7153] = -9'sd187;
	qsin_lut[7154] = -9'sd73;
	icos_lut[7154] = -9'sd176;
	qsin_lut[7155] = -9'sd106;
	icos_lut[7155] = -9'sd159;
	qsin_lut[7156] = -9'sd135;
	icos_lut[7156] = -9'sd135;
	qsin_lut[7157] = -9'sd159;
	icos_lut[7157] = -9'sd106;
	qsin_lut[7158] = -9'sd176;
	icos_lut[7158] = -9'sd73;
	qsin_lut[7159] = -9'sd187;
	icos_lut[7159] = -9'sd37;
	qsin_lut[7160] = -9'sd191;
	icos_lut[7160] = -9'sd0;
	qsin_lut[7161] = -9'sd187;
	icos_lut[7161] =  9'sd37;
	qsin_lut[7162] = -9'sd176;
	icos_lut[7162] =  9'sd73;
	qsin_lut[7163] = -9'sd159;
	icos_lut[7163] =  9'sd106;
	qsin_lut[7164] = -9'sd135;
	icos_lut[7164] =  9'sd135;
	qsin_lut[7165] = -9'sd106;
	icos_lut[7165] =  9'sd159;
	qsin_lut[7166] = -9'sd73;
	icos_lut[7166] =  9'sd176;
	qsin_lut[7167] = -9'sd37;
	icos_lut[7167] =  9'sd187;
	qsin_lut[7168] =  9'sd0;
	icos_lut[7168] =  9'sd193;
	qsin_lut[7169] =  9'sd38;
	icos_lut[7169] =  9'sd189;
	qsin_lut[7170] =  9'sd74;
	icos_lut[7170] =  9'sd178;
	qsin_lut[7171] =  9'sd107;
	icos_lut[7171] =  9'sd160;
	qsin_lut[7172] =  9'sd136;
	icos_lut[7172] =  9'sd136;
	qsin_lut[7173] =  9'sd160;
	icos_lut[7173] =  9'sd107;
	qsin_lut[7174] =  9'sd178;
	icos_lut[7174] =  9'sd74;
	qsin_lut[7175] =  9'sd189;
	icos_lut[7175] =  9'sd38;
	qsin_lut[7176] =  9'sd193;
	icos_lut[7176] =  9'sd0;
	qsin_lut[7177] =  9'sd189;
	icos_lut[7177] = -9'sd38;
	qsin_lut[7178] =  9'sd178;
	icos_lut[7178] = -9'sd74;
	qsin_lut[7179] =  9'sd160;
	icos_lut[7179] = -9'sd107;
	qsin_lut[7180] =  9'sd136;
	icos_lut[7180] = -9'sd136;
	qsin_lut[7181] =  9'sd107;
	icos_lut[7181] = -9'sd160;
	qsin_lut[7182] =  9'sd74;
	icos_lut[7182] = -9'sd178;
	qsin_lut[7183] =  9'sd38;
	icos_lut[7183] = -9'sd189;
	qsin_lut[7184] =  9'sd0;
	icos_lut[7184] = -9'sd193;
	qsin_lut[7185] = -9'sd38;
	icos_lut[7185] = -9'sd189;
	qsin_lut[7186] = -9'sd74;
	icos_lut[7186] = -9'sd178;
	qsin_lut[7187] = -9'sd107;
	icos_lut[7187] = -9'sd160;
	qsin_lut[7188] = -9'sd136;
	icos_lut[7188] = -9'sd136;
	qsin_lut[7189] = -9'sd160;
	icos_lut[7189] = -9'sd107;
	qsin_lut[7190] = -9'sd178;
	icos_lut[7190] = -9'sd74;
	qsin_lut[7191] = -9'sd189;
	icos_lut[7191] = -9'sd38;
	qsin_lut[7192] = -9'sd193;
	icos_lut[7192] = -9'sd0;
	qsin_lut[7193] = -9'sd189;
	icos_lut[7193] =  9'sd38;
	qsin_lut[7194] = -9'sd178;
	icos_lut[7194] =  9'sd74;
	qsin_lut[7195] = -9'sd160;
	icos_lut[7195] =  9'sd107;
	qsin_lut[7196] = -9'sd136;
	icos_lut[7196] =  9'sd136;
	qsin_lut[7197] = -9'sd107;
	icos_lut[7197] =  9'sd160;
	qsin_lut[7198] = -9'sd74;
	icos_lut[7198] =  9'sd178;
	qsin_lut[7199] = -9'sd38;
	icos_lut[7199] =  9'sd189;
	qsin_lut[7200] =  9'sd0;
	icos_lut[7200] =  9'sd195;
	qsin_lut[7201] =  9'sd38;
	icos_lut[7201] =  9'sd191;
	qsin_lut[7202] =  9'sd75;
	icos_lut[7202] =  9'sd180;
	qsin_lut[7203] =  9'sd108;
	icos_lut[7203] =  9'sd162;
	qsin_lut[7204] =  9'sd138;
	icos_lut[7204] =  9'sd138;
	qsin_lut[7205] =  9'sd162;
	icos_lut[7205] =  9'sd108;
	qsin_lut[7206] =  9'sd180;
	icos_lut[7206] =  9'sd75;
	qsin_lut[7207] =  9'sd191;
	icos_lut[7207] =  9'sd38;
	qsin_lut[7208] =  9'sd195;
	icos_lut[7208] =  9'sd0;
	qsin_lut[7209] =  9'sd191;
	icos_lut[7209] = -9'sd38;
	qsin_lut[7210] =  9'sd180;
	icos_lut[7210] = -9'sd75;
	qsin_lut[7211] =  9'sd162;
	icos_lut[7211] = -9'sd108;
	qsin_lut[7212] =  9'sd138;
	icos_lut[7212] = -9'sd138;
	qsin_lut[7213] =  9'sd108;
	icos_lut[7213] = -9'sd162;
	qsin_lut[7214] =  9'sd75;
	icos_lut[7214] = -9'sd180;
	qsin_lut[7215] =  9'sd38;
	icos_lut[7215] = -9'sd191;
	qsin_lut[7216] =  9'sd0;
	icos_lut[7216] = -9'sd195;
	qsin_lut[7217] = -9'sd38;
	icos_lut[7217] = -9'sd191;
	qsin_lut[7218] = -9'sd75;
	icos_lut[7218] = -9'sd180;
	qsin_lut[7219] = -9'sd108;
	icos_lut[7219] = -9'sd162;
	qsin_lut[7220] = -9'sd138;
	icos_lut[7220] = -9'sd138;
	qsin_lut[7221] = -9'sd162;
	icos_lut[7221] = -9'sd108;
	qsin_lut[7222] = -9'sd180;
	icos_lut[7222] = -9'sd75;
	qsin_lut[7223] = -9'sd191;
	icos_lut[7223] = -9'sd38;
	qsin_lut[7224] = -9'sd195;
	icos_lut[7224] = -9'sd0;
	qsin_lut[7225] = -9'sd191;
	icos_lut[7225] =  9'sd38;
	qsin_lut[7226] = -9'sd180;
	icos_lut[7226] =  9'sd75;
	qsin_lut[7227] = -9'sd162;
	icos_lut[7227] =  9'sd108;
	qsin_lut[7228] = -9'sd138;
	icos_lut[7228] =  9'sd138;
	qsin_lut[7229] = -9'sd108;
	icos_lut[7229] =  9'sd162;
	qsin_lut[7230] = -9'sd75;
	icos_lut[7230] =  9'sd180;
	qsin_lut[7231] = -9'sd38;
	icos_lut[7231] =  9'sd191;
	qsin_lut[7232] =  9'sd0;
	icos_lut[7232] =  9'sd197;
	qsin_lut[7233] =  9'sd38;
	icos_lut[7233] =  9'sd193;
	qsin_lut[7234] =  9'sd75;
	icos_lut[7234] =  9'sd182;
	qsin_lut[7235] =  9'sd109;
	icos_lut[7235] =  9'sd164;
	qsin_lut[7236] =  9'sd139;
	icos_lut[7236] =  9'sd139;
	qsin_lut[7237] =  9'sd164;
	icos_lut[7237] =  9'sd109;
	qsin_lut[7238] =  9'sd182;
	icos_lut[7238] =  9'sd75;
	qsin_lut[7239] =  9'sd193;
	icos_lut[7239] =  9'sd38;
	qsin_lut[7240] =  9'sd197;
	icos_lut[7240] =  9'sd0;
	qsin_lut[7241] =  9'sd193;
	icos_lut[7241] = -9'sd38;
	qsin_lut[7242] =  9'sd182;
	icos_lut[7242] = -9'sd75;
	qsin_lut[7243] =  9'sd164;
	icos_lut[7243] = -9'sd109;
	qsin_lut[7244] =  9'sd139;
	icos_lut[7244] = -9'sd139;
	qsin_lut[7245] =  9'sd109;
	icos_lut[7245] = -9'sd164;
	qsin_lut[7246] =  9'sd75;
	icos_lut[7246] = -9'sd182;
	qsin_lut[7247] =  9'sd38;
	icos_lut[7247] = -9'sd193;
	qsin_lut[7248] =  9'sd0;
	icos_lut[7248] = -9'sd197;
	qsin_lut[7249] = -9'sd38;
	icos_lut[7249] = -9'sd193;
	qsin_lut[7250] = -9'sd75;
	icos_lut[7250] = -9'sd182;
	qsin_lut[7251] = -9'sd109;
	icos_lut[7251] = -9'sd164;
	qsin_lut[7252] = -9'sd139;
	icos_lut[7252] = -9'sd139;
	qsin_lut[7253] = -9'sd164;
	icos_lut[7253] = -9'sd109;
	qsin_lut[7254] = -9'sd182;
	icos_lut[7254] = -9'sd75;
	qsin_lut[7255] = -9'sd193;
	icos_lut[7255] = -9'sd38;
	qsin_lut[7256] = -9'sd197;
	icos_lut[7256] = -9'sd0;
	qsin_lut[7257] = -9'sd193;
	icos_lut[7257] =  9'sd38;
	qsin_lut[7258] = -9'sd182;
	icos_lut[7258] =  9'sd75;
	qsin_lut[7259] = -9'sd164;
	icos_lut[7259] =  9'sd109;
	qsin_lut[7260] = -9'sd139;
	icos_lut[7260] =  9'sd139;
	qsin_lut[7261] = -9'sd109;
	icos_lut[7261] =  9'sd164;
	qsin_lut[7262] = -9'sd75;
	icos_lut[7262] =  9'sd182;
	qsin_lut[7263] = -9'sd38;
	icos_lut[7263] =  9'sd193;
	qsin_lut[7264] =  9'sd0;
	icos_lut[7264] =  9'sd199;
	qsin_lut[7265] =  9'sd39;
	icos_lut[7265] =  9'sd195;
	qsin_lut[7266] =  9'sd76;
	icos_lut[7266] =  9'sd184;
	qsin_lut[7267] =  9'sd111;
	icos_lut[7267] =  9'sd165;
	qsin_lut[7268] =  9'sd141;
	icos_lut[7268] =  9'sd141;
	qsin_lut[7269] =  9'sd165;
	icos_lut[7269] =  9'sd111;
	qsin_lut[7270] =  9'sd184;
	icos_lut[7270] =  9'sd76;
	qsin_lut[7271] =  9'sd195;
	icos_lut[7271] =  9'sd39;
	qsin_lut[7272] =  9'sd199;
	icos_lut[7272] =  9'sd0;
	qsin_lut[7273] =  9'sd195;
	icos_lut[7273] = -9'sd39;
	qsin_lut[7274] =  9'sd184;
	icos_lut[7274] = -9'sd76;
	qsin_lut[7275] =  9'sd165;
	icos_lut[7275] = -9'sd111;
	qsin_lut[7276] =  9'sd141;
	icos_lut[7276] = -9'sd141;
	qsin_lut[7277] =  9'sd111;
	icos_lut[7277] = -9'sd165;
	qsin_lut[7278] =  9'sd76;
	icos_lut[7278] = -9'sd184;
	qsin_lut[7279] =  9'sd39;
	icos_lut[7279] = -9'sd195;
	qsin_lut[7280] =  9'sd0;
	icos_lut[7280] = -9'sd199;
	qsin_lut[7281] = -9'sd39;
	icos_lut[7281] = -9'sd195;
	qsin_lut[7282] = -9'sd76;
	icos_lut[7282] = -9'sd184;
	qsin_lut[7283] = -9'sd111;
	icos_lut[7283] = -9'sd165;
	qsin_lut[7284] = -9'sd141;
	icos_lut[7284] = -9'sd141;
	qsin_lut[7285] = -9'sd165;
	icos_lut[7285] = -9'sd111;
	qsin_lut[7286] = -9'sd184;
	icos_lut[7286] = -9'sd76;
	qsin_lut[7287] = -9'sd195;
	icos_lut[7287] = -9'sd39;
	qsin_lut[7288] = -9'sd199;
	icos_lut[7288] = -9'sd0;
	qsin_lut[7289] = -9'sd195;
	icos_lut[7289] =  9'sd39;
	qsin_lut[7290] = -9'sd184;
	icos_lut[7290] =  9'sd76;
	qsin_lut[7291] = -9'sd165;
	icos_lut[7291] =  9'sd111;
	qsin_lut[7292] = -9'sd141;
	icos_lut[7292] =  9'sd141;
	qsin_lut[7293] = -9'sd111;
	icos_lut[7293] =  9'sd165;
	qsin_lut[7294] = -9'sd76;
	icos_lut[7294] =  9'sd184;
	qsin_lut[7295] = -9'sd39;
	icos_lut[7295] =  9'sd195;
	qsin_lut[7296] =  9'sd0;
	icos_lut[7296] =  9'sd201;
	qsin_lut[7297] =  9'sd39;
	icos_lut[7297] =  9'sd197;
	qsin_lut[7298] =  9'sd77;
	icos_lut[7298] =  9'sd186;
	qsin_lut[7299] =  9'sd112;
	icos_lut[7299] =  9'sd167;
	qsin_lut[7300] =  9'sd142;
	icos_lut[7300] =  9'sd142;
	qsin_lut[7301] =  9'sd167;
	icos_lut[7301] =  9'sd112;
	qsin_lut[7302] =  9'sd186;
	icos_lut[7302] =  9'sd77;
	qsin_lut[7303] =  9'sd197;
	icos_lut[7303] =  9'sd39;
	qsin_lut[7304] =  9'sd201;
	icos_lut[7304] =  9'sd0;
	qsin_lut[7305] =  9'sd197;
	icos_lut[7305] = -9'sd39;
	qsin_lut[7306] =  9'sd186;
	icos_lut[7306] = -9'sd77;
	qsin_lut[7307] =  9'sd167;
	icos_lut[7307] = -9'sd112;
	qsin_lut[7308] =  9'sd142;
	icos_lut[7308] = -9'sd142;
	qsin_lut[7309] =  9'sd112;
	icos_lut[7309] = -9'sd167;
	qsin_lut[7310] =  9'sd77;
	icos_lut[7310] = -9'sd186;
	qsin_lut[7311] =  9'sd39;
	icos_lut[7311] = -9'sd197;
	qsin_lut[7312] =  9'sd0;
	icos_lut[7312] = -9'sd201;
	qsin_lut[7313] = -9'sd39;
	icos_lut[7313] = -9'sd197;
	qsin_lut[7314] = -9'sd77;
	icos_lut[7314] = -9'sd186;
	qsin_lut[7315] = -9'sd112;
	icos_lut[7315] = -9'sd167;
	qsin_lut[7316] = -9'sd142;
	icos_lut[7316] = -9'sd142;
	qsin_lut[7317] = -9'sd167;
	icos_lut[7317] = -9'sd112;
	qsin_lut[7318] = -9'sd186;
	icos_lut[7318] = -9'sd77;
	qsin_lut[7319] = -9'sd197;
	icos_lut[7319] = -9'sd39;
	qsin_lut[7320] = -9'sd201;
	icos_lut[7320] = -9'sd0;
	qsin_lut[7321] = -9'sd197;
	icos_lut[7321] =  9'sd39;
	qsin_lut[7322] = -9'sd186;
	icos_lut[7322] =  9'sd77;
	qsin_lut[7323] = -9'sd167;
	icos_lut[7323] =  9'sd112;
	qsin_lut[7324] = -9'sd142;
	icos_lut[7324] =  9'sd142;
	qsin_lut[7325] = -9'sd112;
	icos_lut[7325] =  9'sd167;
	qsin_lut[7326] = -9'sd77;
	icos_lut[7326] =  9'sd186;
	qsin_lut[7327] = -9'sd39;
	icos_lut[7327] =  9'sd197;
	qsin_lut[7328] =  9'sd0;
	icos_lut[7328] =  9'sd203;
	qsin_lut[7329] =  9'sd40;
	icos_lut[7329] =  9'sd199;
	qsin_lut[7330] =  9'sd78;
	icos_lut[7330] =  9'sd188;
	qsin_lut[7331] =  9'sd113;
	icos_lut[7331] =  9'sd169;
	qsin_lut[7332] =  9'sd144;
	icos_lut[7332] =  9'sd144;
	qsin_lut[7333] =  9'sd169;
	icos_lut[7333] =  9'sd113;
	qsin_lut[7334] =  9'sd188;
	icos_lut[7334] =  9'sd78;
	qsin_lut[7335] =  9'sd199;
	icos_lut[7335] =  9'sd40;
	qsin_lut[7336] =  9'sd203;
	icos_lut[7336] =  9'sd0;
	qsin_lut[7337] =  9'sd199;
	icos_lut[7337] = -9'sd40;
	qsin_lut[7338] =  9'sd188;
	icos_lut[7338] = -9'sd78;
	qsin_lut[7339] =  9'sd169;
	icos_lut[7339] = -9'sd113;
	qsin_lut[7340] =  9'sd144;
	icos_lut[7340] = -9'sd144;
	qsin_lut[7341] =  9'sd113;
	icos_lut[7341] = -9'sd169;
	qsin_lut[7342] =  9'sd78;
	icos_lut[7342] = -9'sd188;
	qsin_lut[7343] =  9'sd40;
	icos_lut[7343] = -9'sd199;
	qsin_lut[7344] =  9'sd0;
	icos_lut[7344] = -9'sd203;
	qsin_lut[7345] = -9'sd40;
	icos_lut[7345] = -9'sd199;
	qsin_lut[7346] = -9'sd78;
	icos_lut[7346] = -9'sd188;
	qsin_lut[7347] = -9'sd113;
	icos_lut[7347] = -9'sd169;
	qsin_lut[7348] = -9'sd144;
	icos_lut[7348] = -9'sd144;
	qsin_lut[7349] = -9'sd169;
	icos_lut[7349] = -9'sd113;
	qsin_lut[7350] = -9'sd188;
	icos_lut[7350] = -9'sd78;
	qsin_lut[7351] = -9'sd199;
	icos_lut[7351] = -9'sd40;
	qsin_lut[7352] = -9'sd203;
	icos_lut[7352] = -9'sd0;
	qsin_lut[7353] = -9'sd199;
	icos_lut[7353] =  9'sd40;
	qsin_lut[7354] = -9'sd188;
	icos_lut[7354] =  9'sd78;
	qsin_lut[7355] = -9'sd169;
	icos_lut[7355] =  9'sd113;
	qsin_lut[7356] = -9'sd144;
	icos_lut[7356] =  9'sd144;
	qsin_lut[7357] = -9'sd113;
	icos_lut[7357] =  9'sd169;
	qsin_lut[7358] = -9'sd78;
	icos_lut[7358] =  9'sd188;
	qsin_lut[7359] = -9'sd40;
	icos_lut[7359] =  9'sd199;
	qsin_lut[7360] =  9'sd0;
	icos_lut[7360] =  9'sd205;
	qsin_lut[7361] =  9'sd40;
	icos_lut[7361] =  9'sd201;
	qsin_lut[7362] =  9'sd78;
	icos_lut[7362] =  9'sd189;
	qsin_lut[7363] =  9'sd114;
	icos_lut[7363] =  9'sd170;
	qsin_lut[7364] =  9'sd145;
	icos_lut[7364] =  9'sd145;
	qsin_lut[7365] =  9'sd170;
	icos_lut[7365] =  9'sd114;
	qsin_lut[7366] =  9'sd189;
	icos_lut[7366] =  9'sd78;
	qsin_lut[7367] =  9'sd201;
	icos_lut[7367] =  9'sd40;
	qsin_lut[7368] =  9'sd205;
	icos_lut[7368] =  9'sd0;
	qsin_lut[7369] =  9'sd201;
	icos_lut[7369] = -9'sd40;
	qsin_lut[7370] =  9'sd189;
	icos_lut[7370] = -9'sd78;
	qsin_lut[7371] =  9'sd170;
	icos_lut[7371] = -9'sd114;
	qsin_lut[7372] =  9'sd145;
	icos_lut[7372] = -9'sd145;
	qsin_lut[7373] =  9'sd114;
	icos_lut[7373] = -9'sd170;
	qsin_lut[7374] =  9'sd78;
	icos_lut[7374] = -9'sd189;
	qsin_lut[7375] =  9'sd40;
	icos_lut[7375] = -9'sd201;
	qsin_lut[7376] =  9'sd0;
	icos_lut[7376] = -9'sd205;
	qsin_lut[7377] = -9'sd40;
	icos_lut[7377] = -9'sd201;
	qsin_lut[7378] = -9'sd78;
	icos_lut[7378] = -9'sd189;
	qsin_lut[7379] = -9'sd114;
	icos_lut[7379] = -9'sd170;
	qsin_lut[7380] = -9'sd145;
	icos_lut[7380] = -9'sd145;
	qsin_lut[7381] = -9'sd170;
	icos_lut[7381] = -9'sd114;
	qsin_lut[7382] = -9'sd189;
	icos_lut[7382] = -9'sd78;
	qsin_lut[7383] = -9'sd201;
	icos_lut[7383] = -9'sd40;
	qsin_lut[7384] = -9'sd205;
	icos_lut[7384] = -9'sd0;
	qsin_lut[7385] = -9'sd201;
	icos_lut[7385] =  9'sd40;
	qsin_lut[7386] = -9'sd189;
	icos_lut[7386] =  9'sd78;
	qsin_lut[7387] = -9'sd170;
	icos_lut[7387] =  9'sd114;
	qsin_lut[7388] = -9'sd145;
	icos_lut[7388] =  9'sd145;
	qsin_lut[7389] = -9'sd114;
	icos_lut[7389] =  9'sd170;
	qsin_lut[7390] = -9'sd78;
	icos_lut[7390] =  9'sd189;
	qsin_lut[7391] = -9'sd40;
	icos_lut[7391] =  9'sd201;
	qsin_lut[7392] =  9'sd0;
	icos_lut[7392] =  9'sd207;
	qsin_lut[7393] =  9'sd40;
	icos_lut[7393] =  9'sd203;
	qsin_lut[7394] =  9'sd79;
	icos_lut[7394] =  9'sd191;
	qsin_lut[7395] =  9'sd115;
	icos_lut[7395] =  9'sd172;
	qsin_lut[7396] =  9'sd146;
	icos_lut[7396] =  9'sd146;
	qsin_lut[7397] =  9'sd172;
	icos_lut[7397] =  9'sd115;
	qsin_lut[7398] =  9'sd191;
	icos_lut[7398] =  9'sd79;
	qsin_lut[7399] =  9'sd203;
	icos_lut[7399] =  9'sd40;
	qsin_lut[7400] =  9'sd207;
	icos_lut[7400] =  9'sd0;
	qsin_lut[7401] =  9'sd203;
	icos_lut[7401] = -9'sd40;
	qsin_lut[7402] =  9'sd191;
	icos_lut[7402] = -9'sd79;
	qsin_lut[7403] =  9'sd172;
	icos_lut[7403] = -9'sd115;
	qsin_lut[7404] =  9'sd146;
	icos_lut[7404] = -9'sd146;
	qsin_lut[7405] =  9'sd115;
	icos_lut[7405] = -9'sd172;
	qsin_lut[7406] =  9'sd79;
	icos_lut[7406] = -9'sd191;
	qsin_lut[7407] =  9'sd40;
	icos_lut[7407] = -9'sd203;
	qsin_lut[7408] =  9'sd0;
	icos_lut[7408] = -9'sd207;
	qsin_lut[7409] = -9'sd40;
	icos_lut[7409] = -9'sd203;
	qsin_lut[7410] = -9'sd79;
	icos_lut[7410] = -9'sd191;
	qsin_lut[7411] = -9'sd115;
	icos_lut[7411] = -9'sd172;
	qsin_lut[7412] = -9'sd146;
	icos_lut[7412] = -9'sd146;
	qsin_lut[7413] = -9'sd172;
	icos_lut[7413] = -9'sd115;
	qsin_lut[7414] = -9'sd191;
	icos_lut[7414] = -9'sd79;
	qsin_lut[7415] = -9'sd203;
	icos_lut[7415] = -9'sd40;
	qsin_lut[7416] = -9'sd207;
	icos_lut[7416] = -9'sd0;
	qsin_lut[7417] = -9'sd203;
	icos_lut[7417] =  9'sd40;
	qsin_lut[7418] = -9'sd191;
	icos_lut[7418] =  9'sd79;
	qsin_lut[7419] = -9'sd172;
	icos_lut[7419] =  9'sd115;
	qsin_lut[7420] = -9'sd146;
	icos_lut[7420] =  9'sd146;
	qsin_lut[7421] = -9'sd115;
	icos_lut[7421] =  9'sd172;
	qsin_lut[7422] = -9'sd79;
	icos_lut[7422] =  9'sd191;
	qsin_lut[7423] = -9'sd40;
	icos_lut[7423] =  9'sd203;
	qsin_lut[7424] =  9'sd0;
	icos_lut[7424] =  9'sd209;
	qsin_lut[7425] =  9'sd41;
	icos_lut[7425] =  9'sd205;
	qsin_lut[7426] =  9'sd80;
	icos_lut[7426] =  9'sd193;
	qsin_lut[7427] =  9'sd116;
	icos_lut[7427] =  9'sd174;
	qsin_lut[7428] =  9'sd148;
	icos_lut[7428] =  9'sd148;
	qsin_lut[7429] =  9'sd174;
	icos_lut[7429] =  9'sd116;
	qsin_lut[7430] =  9'sd193;
	icos_lut[7430] =  9'sd80;
	qsin_lut[7431] =  9'sd205;
	icos_lut[7431] =  9'sd41;
	qsin_lut[7432] =  9'sd209;
	icos_lut[7432] =  9'sd0;
	qsin_lut[7433] =  9'sd205;
	icos_lut[7433] = -9'sd41;
	qsin_lut[7434] =  9'sd193;
	icos_lut[7434] = -9'sd80;
	qsin_lut[7435] =  9'sd174;
	icos_lut[7435] = -9'sd116;
	qsin_lut[7436] =  9'sd148;
	icos_lut[7436] = -9'sd148;
	qsin_lut[7437] =  9'sd116;
	icos_lut[7437] = -9'sd174;
	qsin_lut[7438] =  9'sd80;
	icos_lut[7438] = -9'sd193;
	qsin_lut[7439] =  9'sd41;
	icos_lut[7439] = -9'sd205;
	qsin_lut[7440] =  9'sd0;
	icos_lut[7440] = -9'sd209;
	qsin_lut[7441] = -9'sd41;
	icos_lut[7441] = -9'sd205;
	qsin_lut[7442] = -9'sd80;
	icos_lut[7442] = -9'sd193;
	qsin_lut[7443] = -9'sd116;
	icos_lut[7443] = -9'sd174;
	qsin_lut[7444] = -9'sd148;
	icos_lut[7444] = -9'sd148;
	qsin_lut[7445] = -9'sd174;
	icos_lut[7445] = -9'sd116;
	qsin_lut[7446] = -9'sd193;
	icos_lut[7446] = -9'sd80;
	qsin_lut[7447] = -9'sd205;
	icos_lut[7447] = -9'sd41;
	qsin_lut[7448] = -9'sd209;
	icos_lut[7448] = -9'sd0;
	qsin_lut[7449] = -9'sd205;
	icos_lut[7449] =  9'sd41;
	qsin_lut[7450] = -9'sd193;
	icos_lut[7450] =  9'sd80;
	qsin_lut[7451] = -9'sd174;
	icos_lut[7451] =  9'sd116;
	qsin_lut[7452] = -9'sd148;
	icos_lut[7452] =  9'sd148;
	qsin_lut[7453] = -9'sd116;
	icos_lut[7453] =  9'sd174;
	qsin_lut[7454] = -9'sd80;
	icos_lut[7454] =  9'sd193;
	qsin_lut[7455] = -9'sd41;
	icos_lut[7455] =  9'sd205;
	qsin_lut[7456] =  9'sd0;
	icos_lut[7456] =  9'sd211;
	qsin_lut[7457] =  9'sd41;
	icos_lut[7457] =  9'sd207;
	qsin_lut[7458] =  9'sd81;
	icos_lut[7458] =  9'sd195;
	qsin_lut[7459] =  9'sd117;
	icos_lut[7459] =  9'sd175;
	qsin_lut[7460] =  9'sd149;
	icos_lut[7460] =  9'sd149;
	qsin_lut[7461] =  9'sd175;
	icos_lut[7461] =  9'sd117;
	qsin_lut[7462] =  9'sd195;
	icos_lut[7462] =  9'sd81;
	qsin_lut[7463] =  9'sd207;
	icos_lut[7463] =  9'sd41;
	qsin_lut[7464] =  9'sd211;
	icos_lut[7464] =  9'sd0;
	qsin_lut[7465] =  9'sd207;
	icos_lut[7465] = -9'sd41;
	qsin_lut[7466] =  9'sd195;
	icos_lut[7466] = -9'sd81;
	qsin_lut[7467] =  9'sd175;
	icos_lut[7467] = -9'sd117;
	qsin_lut[7468] =  9'sd149;
	icos_lut[7468] = -9'sd149;
	qsin_lut[7469] =  9'sd117;
	icos_lut[7469] = -9'sd175;
	qsin_lut[7470] =  9'sd81;
	icos_lut[7470] = -9'sd195;
	qsin_lut[7471] =  9'sd41;
	icos_lut[7471] = -9'sd207;
	qsin_lut[7472] =  9'sd0;
	icos_lut[7472] = -9'sd211;
	qsin_lut[7473] = -9'sd41;
	icos_lut[7473] = -9'sd207;
	qsin_lut[7474] = -9'sd81;
	icos_lut[7474] = -9'sd195;
	qsin_lut[7475] = -9'sd117;
	icos_lut[7475] = -9'sd175;
	qsin_lut[7476] = -9'sd149;
	icos_lut[7476] = -9'sd149;
	qsin_lut[7477] = -9'sd175;
	icos_lut[7477] = -9'sd117;
	qsin_lut[7478] = -9'sd195;
	icos_lut[7478] = -9'sd81;
	qsin_lut[7479] = -9'sd207;
	icos_lut[7479] = -9'sd41;
	qsin_lut[7480] = -9'sd211;
	icos_lut[7480] = -9'sd0;
	qsin_lut[7481] = -9'sd207;
	icos_lut[7481] =  9'sd41;
	qsin_lut[7482] = -9'sd195;
	icos_lut[7482] =  9'sd81;
	qsin_lut[7483] = -9'sd175;
	icos_lut[7483] =  9'sd117;
	qsin_lut[7484] = -9'sd149;
	icos_lut[7484] =  9'sd149;
	qsin_lut[7485] = -9'sd117;
	icos_lut[7485] =  9'sd175;
	qsin_lut[7486] = -9'sd81;
	icos_lut[7486] =  9'sd195;
	qsin_lut[7487] = -9'sd41;
	icos_lut[7487] =  9'sd207;
	qsin_lut[7488] =  9'sd0;
	icos_lut[7488] =  9'sd213;
	qsin_lut[7489] =  9'sd42;
	icos_lut[7489] =  9'sd209;
	qsin_lut[7490] =  9'sd82;
	icos_lut[7490] =  9'sd197;
	qsin_lut[7491] =  9'sd118;
	icos_lut[7491] =  9'sd177;
	qsin_lut[7492] =  9'sd151;
	icos_lut[7492] =  9'sd151;
	qsin_lut[7493] =  9'sd177;
	icos_lut[7493] =  9'sd118;
	qsin_lut[7494] =  9'sd197;
	icos_lut[7494] =  9'sd82;
	qsin_lut[7495] =  9'sd209;
	icos_lut[7495] =  9'sd42;
	qsin_lut[7496] =  9'sd213;
	icos_lut[7496] =  9'sd0;
	qsin_lut[7497] =  9'sd209;
	icos_lut[7497] = -9'sd42;
	qsin_lut[7498] =  9'sd197;
	icos_lut[7498] = -9'sd82;
	qsin_lut[7499] =  9'sd177;
	icos_lut[7499] = -9'sd118;
	qsin_lut[7500] =  9'sd151;
	icos_lut[7500] = -9'sd151;
	qsin_lut[7501] =  9'sd118;
	icos_lut[7501] = -9'sd177;
	qsin_lut[7502] =  9'sd82;
	icos_lut[7502] = -9'sd197;
	qsin_lut[7503] =  9'sd42;
	icos_lut[7503] = -9'sd209;
	qsin_lut[7504] =  9'sd0;
	icos_lut[7504] = -9'sd213;
	qsin_lut[7505] = -9'sd42;
	icos_lut[7505] = -9'sd209;
	qsin_lut[7506] = -9'sd82;
	icos_lut[7506] = -9'sd197;
	qsin_lut[7507] = -9'sd118;
	icos_lut[7507] = -9'sd177;
	qsin_lut[7508] = -9'sd151;
	icos_lut[7508] = -9'sd151;
	qsin_lut[7509] = -9'sd177;
	icos_lut[7509] = -9'sd118;
	qsin_lut[7510] = -9'sd197;
	icos_lut[7510] = -9'sd82;
	qsin_lut[7511] = -9'sd209;
	icos_lut[7511] = -9'sd42;
	qsin_lut[7512] = -9'sd213;
	icos_lut[7512] = -9'sd0;
	qsin_lut[7513] = -9'sd209;
	icos_lut[7513] =  9'sd42;
	qsin_lut[7514] = -9'sd197;
	icos_lut[7514] =  9'sd82;
	qsin_lut[7515] = -9'sd177;
	icos_lut[7515] =  9'sd118;
	qsin_lut[7516] = -9'sd151;
	icos_lut[7516] =  9'sd151;
	qsin_lut[7517] = -9'sd118;
	icos_lut[7517] =  9'sd177;
	qsin_lut[7518] = -9'sd82;
	icos_lut[7518] =  9'sd197;
	qsin_lut[7519] = -9'sd42;
	icos_lut[7519] =  9'sd209;
	qsin_lut[7520] =  9'sd0;
	icos_lut[7520] =  9'sd215;
	qsin_lut[7521] =  9'sd42;
	icos_lut[7521] =  9'sd211;
	qsin_lut[7522] =  9'sd82;
	icos_lut[7522] =  9'sd199;
	qsin_lut[7523] =  9'sd119;
	icos_lut[7523] =  9'sd179;
	qsin_lut[7524] =  9'sd152;
	icos_lut[7524] =  9'sd152;
	qsin_lut[7525] =  9'sd179;
	icos_lut[7525] =  9'sd119;
	qsin_lut[7526] =  9'sd199;
	icos_lut[7526] =  9'sd82;
	qsin_lut[7527] =  9'sd211;
	icos_lut[7527] =  9'sd42;
	qsin_lut[7528] =  9'sd215;
	icos_lut[7528] =  9'sd0;
	qsin_lut[7529] =  9'sd211;
	icos_lut[7529] = -9'sd42;
	qsin_lut[7530] =  9'sd199;
	icos_lut[7530] = -9'sd82;
	qsin_lut[7531] =  9'sd179;
	icos_lut[7531] = -9'sd119;
	qsin_lut[7532] =  9'sd152;
	icos_lut[7532] = -9'sd152;
	qsin_lut[7533] =  9'sd119;
	icos_lut[7533] = -9'sd179;
	qsin_lut[7534] =  9'sd82;
	icos_lut[7534] = -9'sd199;
	qsin_lut[7535] =  9'sd42;
	icos_lut[7535] = -9'sd211;
	qsin_lut[7536] =  9'sd0;
	icos_lut[7536] = -9'sd215;
	qsin_lut[7537] = -9'sd42;
	icos_lut[7537] = -9'sd211;
	qsin_lut[7538] = -9'sd82;
	icos_lut[7538] = -9'sd199;
	qsin_lut[7539] = -9'sd119;
	icos_lut[7539] = -9'sd179;
	qsin_lut[7540] = -9'sd152;
	icos_lut[7540] = -9'sd152;
	qsin_lut[7541] = -9'sd179;
	icos_lut[7541] = -9'sd119;
	qsin_lut[7542] = -9'sd199;
	icos_lut[7542] = -9'sd82;
	qsin_lut[7543] = -9'sd211;
	icos_lut[7543] = -9'sd42;
	qsin_lut[7544] = -9'sd215;
	icos_lut[7544] = -9'sd0;
	qsin_lut[7545] = -9'sd211;
	icos_lut[7545] =  9'sd42;
	qsin_lut[7546] = -9'sd199;
	icos_lut[7546] =  9'sd82;
	qsin_lut[7547] = -9'sd179;
	icos_lut[7547] =  9'sd119;
	qsin_lut[7548] = -9'sd152;
	icos_lut[7548] =  9'sd152;
	qsin_lut[7549] = -9'sd119;
	icos_lut[7549] =  9'sd179;
	qsin_lut[7550] = -9'sd82;
	icos_lut[7550] =  9'sd199;
	qsin_lut[7551] = -9'sd42;
	icos_lut[7551] =  9'sd211;
	qsin_lut[7552] =  9'sd0;
	icos_lut[7552] =  9'sd217;
	qsin_lut[7553] =  9'sd42;
	icos_lut[7553] =  9'sd213;
	qsin_lut[7554] =  9'sd83;
	icos_lut[7554] =  9'sd200;
	qsin_lut[7555] =  9'sd121;
	icos_lut[7555] =  9'sd180;
	qsin_lut[7556] =  9'sd153;
	icos_lut[7556] =  9'sd153;
	qsin_lut[7557] =  9'sd180;
	icos_lut[7557] =  9'sd121;
	qsin_lut[7558] =  9'sd200;
	icos_lut[7558] =  9'sd83;
	qsin_lut[7559] =  9'sd213;
	icos_lut[7559] =  9'sd42;
	qsin_lut[7560] =  9'sd217;
	icos_lut[7560] =  9'sd0;
	qsin_lut[7561] =  9'sd213;
	icos_lut[7561] = -9'sd42;
	qsin_lut[7562] =  9'sd200;
	icos_lut[7562] = -9'sd83;
	qsin_lut[7563] =  9'sd180;
	icos_lut[7563] = -9'sd121;
	qsin_lut[7564] =  9'sd153;
	icos_lut[7564] = -9'sd153;
	qsin_lut[7565] =  9'sd121;
	icos_lut[7565] = -9'sd180;
	qsin_lut[7566] =  9'sd83;
	icos_lut[7566] = -9'sd200;
	qsin_lut[7567] =  9'sd42;
	icos_lut[7567] = -9'sd213;
	qsin_lut[7568] =  9'sd0;
	icos_lut[7568] = -9'sd217;
	qsin_lut[7569] = -9'sd42;
	icos_lut[7569] = -9'sd213;
	qsin_lut[7570] = -9'sd83;
	icos_lut[7570] = -9'sd200;
	qsin_lut[7571] = -9'sd121;
	icos_lut[7571] = -9'sd180;
	qsin_lut[7572] = -9'sd153;
	icos_lut[7572] = -9'sd153;
	qsin_lut[7573] = -9'sd180;
	icos_lut[7573] = -9'sd121;
	qsin_lut[7574] = -9'sd200;
	icos_lut[7574] = -9'sd83;
	qsin_lut[7575] = -9'sd213;
	icos_lut[7575] = -9'sd42;
	qsin_lut[7576] = -9'sd217;
	icos_lut[7576] = -9'sd0;
	qsin_lut[7577] = -9'sd213;
	icos_lut[7577] =  9'sd42;
	qsin_lut[7578] = -9'sd200;
	icos_lut[7578] =  9'sd83;
	qsin_lut[7579] = -9'sd180;
	icos_lut[7579] =  9'sd121;
	qsin_lut[7580] = -9'sd153;
	icos_lut[7580] =  9'sd153;
	qsin_lut[7581] = -9'sd121;
	icos_lut[7581] =  9'sd180;
	qsin_lut[7582] = -9'sd83;
	icos_lut[7582] =  9'sd200;
	qsin_lut[7583] = -9'sd42;
	icos_lut[7583] =  9'sd213;
	qsin_lut[7584] =  9'sd0;
	icos_lut[7584] =  9'sd219;
	qsin_lut[7585] =  9'sd43;
	icos_lut[7585] =  9'sd215;
	qsin_lut[7586] =  9'sd84;
	icos_lut[7586] =  9'sd202;
	qsin_lut[7587] =  9'sd122;
	icos_lut[7587] =  9'sd182;
	qsin_lut[7588] =  9'sd155;
	icos_lut[7588] =  9'sd155;
	qsin_lut[7589] =  9'sd182;
	icos_lut[7589] =  9'sd122;
	qsin_lut[7590] =  9'sd202;
	icos_lut[7590] =  9'sd84;
	qsin_lut[7591] =  9'sd215;
	icos_lut[7591] =  9'sd43;
	qsin_lut[7592] =  9'sd219;
	icos_lut[7592] =  9'sd0;
	qsin_lut[7593] =  9'sd215;
	icos_lut[7593] = -9'sd43;
	qsin_lut[7594] =  9'sd202;
	icos_lut[7594] = -9'sd84;
	qsin_lut[7595] =  9'sd182;
	icos_lut[7595] = -9'sd122;
	qsin_lut[7596] =  9'sd155;
	icos_lut[7596] = -9'sd155;
	qsin_lut[7597] =  9'sd122;
	icos_lut[7597] = -9'sd182;
	qsin_lut[7598] =  9'sd84;
	icos_lut[7598] = -9'sd202;
	qsin_lut[7599] =  9'sd43;
	icos_lut[7599] = -9'sd215;
	qsin_lut[7600] =  9'sd0;
	icos_lut[7600] = -9'sd219;
	qsin_lut[7601] = -9'sd43;
	icos_lut[7601] = -9'sd215;
	qsin_lut[7602] = -9'sd84;
	icos_lut[7602] = -9'sd202;
	qsin_lut[7603] = -9'sd122;
	icos_lut[7603] = -9'sd182;
	qsin_lut[7604] = -9'sd155;
	icos_lut[7604] = -9'sd155;
	qsin_lut[7605] = -9'sd182;
	icos_lut[7605] = -9'sd122;
	qsin_lut[7606] = -9'sd202;
	icos_lut[7606] = -9'sd84;
	qsin_lut[7607] = -9'sd215;
	icos_lut[7607] = -9'sd43;
	qsin_lut[7608] = -9'sd219;
	icos_lut[7608] = -9'sd0;
	qsin_lut[7609] = -9'sd215;
	icos_lut[7609] =  9'sd43;
	qsin_lut[7610] = -9'sd202;
	icos_lut[7610] =  9'sd84;
	qsin_lut[7611] = -9'sd182;
	icos_lut[7611] =  9'sd122;
	qsin_lut[7612] = -9'sd155;
	icos_lut[7612] =  9'sd155;
	qsin_lut[7613] = -9'sd122;
	icos_lut[7613] =  9'sd182;
	qsin_lut[7614] = -9'sd84;
	icos_lut[7614] =  9'sd202;
	qsin_lut[7615] = -9'sd43;
	icos_lut[7615] =  9'sd215;
	qsin_lut[7616] =  9'sd0;
	icos_lut[7616] =  9'sd221;
	qsin_lut[7617] =  9'sd43;
	icos_lut[7617] =  9'sd217;
	qsin_lut[7618] =  9'sd85;
	icos_lut[7618] =  9'sd204;
	qsin_lut[7619] =  9'sd123;
	icos_lut[7619] =  9'sd184;
	qsin_lut[7620] =  9'sd156;
	icos_lut[7620] =  9'sd156;
	qsin_lut[7621] =  9'sd184;
	icos_lut[7621] =  9'sd123;
	qsin_lut[7622] =  9'sd204;
	icos_lut[7622] =  9'sd85;
	qsin_lut[7623] =  9'sd217;
	icos_lut[7623] =  9'sd43;
	qsin_lut[7624] =  9'sd221;
	icos_lut[7624] =  9'sd0;
	qsin_lut[7625] =  9'sd217;
	icos_lut[7625] = -9'sd43;
	qsin_lut[7626] =  9'sd204;
	icos_lut[7626] = -9'sd85;
	qsin_lut[7627] =  9'sd184;
	icos_lut[7627] = -9'sd123;
	qsin_lut[7628] =  9'sd156;
	icos_lut[7628] = -9'sd156;
	qsin_lut[7629] =  9'sd123;
	icos_lut[7629] = -9'sd184;
	qsin_lut[7630] =  9'sd85;
	icos_lut[7630] = -9'sd204;
	qsin_lut[7631] =  9'sd43;
	icos_lut[7631] = -9'sd217;
	qsin_lut[7632] =  9'sd0;
	icos_lut[7632] = -9'sd221;
	qsin_lut[7633] = -9'sd43;
	icos_lut[7633] = -9'sd217;
	qsin_lut[7634] = -9'sd85;
	icos_lut[7634] = -9'sd204;
	qsin_lut[7635] = -9'sd123;
	icos_lut[7635] = -9'sd184;
	qsin_lut[7636] = -9'sd156;
	icos_lut[7636] = -9'sd156;
	qsin_lut[7637] = -9'sd184;
	icos_lut[7637] = -9'sd123;
	qsin_lut[7638] = -9'sd204;
	icos_lut[7638] = -9'sd85;
	qsin_lut[7639] = -9'sd217;
	icos_lut[7639] = -9'sd43;
	qsin_lut[7640] = -9'sd221;
	icos_lut[7640] = -9'sd0;
	qsin_lut[7641] = -9'sd217;
	icos_lut[7641] =  9'sd43;
	qsin_lut[7642] = -9'sd204;
	icos_lut[7642] =  9'sd85;
	qsin_lut[7643] = -9'sd184;
	icos_lut[7643] =  9'sd123;
	qsin_lut[7644] = -9'sd156;
	icos_lut[7644] =  9'sd156;
	qsin_lut[7645] = -9'sd123;
	icos_lut[7645] =  9'sd184;
	qsin_lut[7646] = -9'sd85;
	icos_lut[7646] =  9'sd204;
	qsin_lut[7647] = -9'sd43;
	icos_lut[7647] =  9'sd217;
	qsin_lut[7648] =  9'sd0;
	icos_lut[7648] =  9'sd223;
	qsin_lut[7649] =  9'sd44;
	icos_lut[7649] =  9'sd219;
	qsin_lut[7650] =  9'sd85;
	icos_lut[7650] =  9'sd206;
	qsin_lut[7651] =  9'sd124;
	icos_lut[7651] =  9'sd185;
	qsin_lut[7652] =  9'sd158;
	icos_lut[7652] =  9'sd158;
	qsin_lut[7653] =  9'sd185;
	icos_lut[7653] =  9'sd124;
	qsin_lut[7654] =  9'sd206;
	icos_lut[7654] =  9'sd85;
	qsin_lut[7655] =  9'sd219;
	icos_lut[7655] =  9'sd44;
	qsin_lut[7656] =  9'sd223;
	icos_lut[7656] =  9'sd0;
	qsin_lut[7657] =  9'sd219;
	icos_lut[7657] = -9'sd44;
	qsin_lut[7658] =  9'sd206;
	icos_lut[7658] = -9'sd85;
	qsin_lut[7659] =  9'sd185;
	icos_lut[7659] = -9'sd124;
	qsin_lut[7660] =  9'sd158;
	icos_lut[7660] = -9'sd158;
	qsin_lut[7661] =  9'sd124;
	icos_lut[7661] = -9'sd185;
	qsin_lut[7662] =  9'sd85;
	icos_lut[7662] = -9'sd206;
	qsin_lut[7663] =  9'sd44;
	icos_lut[7663] = -9'sd219;
	qsin_lut[7664] =  9'sd0;
	icos_lut[7664] = -9'sd223;
	qsin_lut[7665] = -9'sd44;
	icos_lut[7665] = -9'sd219;
	qsin_lut[7666] = -9'sd85;
	icos_lut[7666] = -9'sd206;
	qsin_lut[7667] = -9'sd124;
	icos_lut[7667] = -9'sd185;
	qsin_lut[7668] = -9'sd158;
	icos_lut[7668] = -9'sd158;
	qsin_lut[7669] = -9'sd185;
	icos_lut[7669] = -9'sd124;
	qsin_lut[7670] = -9'sd206;
	icos_lut[7670] = -9'sd85;
	qsin_lut[7671] = -9'sd219;
	icos_lut[7671] = -9'sd44;
	qsin_lut[7672] = -9'sd223;
	icos_lut[7672] = -9'sd0;
	qsin_lut[7673] = -9'sd219;
	icos_lut[7673] =  9'sd44;
	qsin_lut[7674] = -9'sd206;
	icos_lut[7674] =  9'sd85;
	qsin_lut[7675] = -9'sd185;
	icos_lut[7675] =  9'sd124;
	qsin_lut[7676] = -9'sd158;
	icos_lut[7676] =  9'sd158;
	qsin_lut[7677] = -9'sd124;
	icos_lut[7677] =  9'sd185;
	qsin_lut[7678] = -9'sd85;
	icos_lut[7678] =  9'sd206;
	qsin_lut[7679] = -9'sd44;
	icos_lut[7679] =  9'sd219;
	qsin_lut[7680] =  9'sd0;
	icos_lut[7680] =  9'sd225;
	qsin_lut[7681] =  9'sd44;
	icos_lut[7681] =  9'sd221;
	qsin_lut[7682] =  9'sd86;
	icos_lut[7682] =  9'sd208;
	qsin_lut[7683] =  9'sd125;
	icos_lut[7683] =  9'sd187;
	qsin_lut[7684] =  9'sd159;
	icos_lut[7684] =  9'sd159;
	qsin_lut[7685] =  9'sd187;
	icos_lut[7685] =  9'sd125;
	qsin_lut[7686] =  9'sd208;
	icos_lut[7686] =  9'sd86;
	qsin_lut[7687] =  9'sd221;
	icos_lut[7687] =  9'sd44;
	qsin_lut[7688] =  9'sd225;
	icos_lut[7688] =  9'sd0;
	qsin_lut[7689] =  9'sd221;
	icos_lut[7689] = -9'sd44;
	qsin_lut[7690] =  9'sd208;
	icos_lut[7690] = -9'sd86;
	qsin_lut[7691] =  9'sd187;
	icos_lut[7691] = -9'sd125;
	qsin_lut[7692] =  9'sd159;
	icos_lut[7692] = -9'sd159;
	qsin_lut[7693] =  9'sd125;
	icos_lut[7693] = -9'sd187;
	qsin_lut[7694] =  9'sd86;
	icos_lut[7694] = -9'sd208;
	qsin_lut[7695] =  9'sd44;
	icos_lut[7695] = -9'sd221;
	qsin_lut[7696] =  9'sd0;
	icos_lut[7696] = -9'sd225;
	qsin_lut[7697] = -9'sd44;
	icos_lut[7697] = -9'sd221;
	qsin_lut[7698] = -9'sd86;
	icos_lut[7698] = -9'sd208;
	qsin_lut[7699] = -9'sd125;
	icos_lut[7699] = -9'sd187;
	qsin_lut[7700] = -9'sd159;
	icos_lut[7700] = -9'sd159;
	qsin_lut[7701] = -9'sd187;
	icos_lut[7701] = -9'sd125;
	qsin_lut[7702] = -9'sd208;
	icos_lut[7702] = -9'sd86;
	qsin_lut[7703] = -9'sd221;
	icos_lut[7703] = -9'sd44;
	qsin_lut[7704] = -9'sd225;
	icos_lut[7704] = -9'sd0;
	qsin_lut[7705] = -9'sd221;
	icos_lut[7705] =  9'sd44;
	qsin_lut[7706] = -9'sd208;
	icos_lut[7706] =  9'sd86;
	qsin_lut[7707] = -9'sd187;
	icos_lut[7707] =  9'sd125;
	qsin_lut[7708] = -9'sd159;
	icos_lut[7708] =  9'sd159;
	qsin_lut[7709] = -9'sd125;
	icos_lut[7709] =  9'sd187;
	qsin_lut[7710] = -9'sd86;
	icos_lut[7710] =  9'sd208;
	qsin_lut[7711] = -9'sd44;
	icos_lut[7711] =  9'sd221;
	qsin_lut[7712] =  9'sd0;
	icos_lut[7712] =  9'sd227;
	qsin_lut[7713] =  9'sd44;
	icos_lut[7713] =  9'sd223;
	qsin_lut[7714] =  9'sd87;
	icos_lut[7714] =  9'sd210;
	qsin_lut[7715] =  9'sd126;
	icos_lut[7715] =  9'sd189;
	qsin_lut[7716] =  9'sd161;
	icos_lut[7716] =  9'sd161;
	qsin_lut[7717] =  9'sd189;
	icos_lut[7717] =  9'sd126;
	qsin_lut[7718] =  9'sd210;
	icos_lut[7718] =  9'sd87;
	qsin_lut[7719] =  9'sd223;
	icos_lut[7719] =  9'sd44;
	qsin_lut[7720] =  9'sd227;
	icos_lut[7720] =  9'sd0;
	qsin_lut[7721] =  9'sd223;
	icos_lut[7721] = -9'sd44;
	qsin_lut[7722] =  9'sd210;
	icos_lut[7722] = -9'sd87;
	qsin_lut[7723] =  9'sd189;
	icos_lut[7723] = -9'sd126;
	qsin_lut[7724] =  9'sd161;
	icos_lut[7724] = -9'sd161;
	qsin_lut[7725] =  9'sd126;
	icos_lut[7725] = -9'sd189;
	qsin_lut[7726] =  9'sd87;
	icos_lut[7726] = -9'sd210;
	qsin_lut[7727] =  9'sd44;
	icos_lut[7727] = -9'sd223;
	qsin_lut[7728] =  9'sd0;
	icos_lut[7728] = -9'sd227;
	qsin_lut[7729] = -9'sd44;
	icos_lut[7729] = -9'sd223;
	qsin_lut[7730] = -9'sd87;
	icos_lut[7730] = -9'sd210;
	qsin_lut[7731] = -9'sd126;
	icos_lut[7731] = -9'sd189;
	qsin_lut[7732] = -9'sd161;
	icos_lut[7732] = -9'sd161;
	qsin_lut[7733] = -9'sd189;
	icos_lut[7733] = -9'sd126;
	qsin_lut[7734] = -9'sd210;
	icos_lut[7734] = -9'sd87;
	qsin_lut[7735] = -9'sd223;
	icos_lut[7735] = -9'sd44;
	qsin_lut[7736] = -9'sd227;
	icos_lut[7736] = -9'sd0;
	qsin_lut[7737] = -9'sd223;
	icos_lut[7737] =  9'sd44;
	qsin_lut[7738] = -9'sd210;
	icos_lut[7738] =  9'sd87;
	qsin_lut[7739] = -9'sd189;
	icos_lut[7739] =  9'sd126;
	qsin_lut[7740] = -9'sd161;
	icos_lut[7740] =  9'sd161;
	qsin_lut[7741] = -9'sd126;
	icos_lut[7741] =  9'sd189;
	qsin_lut[7742] = -9'sd87;
	icos_lut[7742] =  9'sd210;
	qsin_lut[7743] = -9'sd44;
	icos_lut[7743] =  9'sd223;
	qsin_lut[7744] =  9'sd0;
	icos_lut[7744] =  9'sd229;
	qsin_lut[7745] =  9'sd45;
	icos_lut[7745] =  9'sd225;
	qsin_lut[7746] =  9'sd88;
	icos_lut[7746] =  9'sd212;
	qsin_lut[7747] =  9'sd127;
	icos_lut[7747] =  9'sd190;
	qsin_lut[7748] =  9'sd162;
	icos_lut[7748] =  9'sd162;
	qsin_lut[7749] =  9'sd190;
	icos_lut[7749] =  9'sd127;
	qsin_lut[7750] =  9'sd212;
	icos_lut[7750] =  9'sd88;
	qsin_lut[7751] =  9'sd225;
	icos_lut[7751] =  9'sd45;
	qsin_lut[7752] =  9'sd229;
	icos_lut[7752] =  9'sd0;
	qsin_lut[7753] =  9'sd225;
	icos_lut[7753] = -9'sd45;
	qsin_lut[7754] =  9'sd212;
	icos_lut[7754] = -9'sd88;
	qsin_lut[7755] =  9'sd190;
	icos_lut[7755] = -9'sd127;
	qsin_lut[7756] =  9'sd162;
	icos_lut[7756] = -9'sd162;
	qsin_lut[7757] =  9'sd127;
	icos_lut[7757] = -9'sd190;
	qsin_lut[7758] =  9'sd88;
	icos_lut[7758] = -9'sd212;
	qsin_lut[7759] =  9'sd45;
	icos_lut[7759] = -9'sd225;
	qsin_lut[7760] =  9'sd0;
	icos_lut[7760] = -9'sd229;
	qsin_lut[7761] = -9'sd45;
	icos_lut[7761] = -9'sd225;
	qsin_lut[7762] = -9'sd88;
	icos_lut[7762] = -9'sd212;
	qsin_lut[7763] = -9'sd127;
	icos_lut[7763] = -9'sd190;
	qsin_lut[7764] = -9'sd162;
	icos_lut[7764] = -9'sd162;
	qsin_lut[7765] = -9'sd190;
	icos_lut[7765] = -9'sd127;
	qsin_lut[7766] = -9'sd212;
	icos_lut[7766] = -9'sd88;
	qsin_lut[7767] = -9'sd225;
	icos_lut[7767] = -9'sd45;
	qsin_lut[7768] = -9'sd229;
	icos_lut[7768] = -9'sd0;
	qsin_lut[7769] = -9'sd225;
	icos_lut[7769] =  9'sd45;
	qsin_lut[7770] = -9'sd212;
	icos_lut[7770] =  9'sd88;
	qsin_lut[7771] = -9'sd190;
	icos_lut[7771] =  9'sd127;
	qsin_lut[7772] = -9'sd162;
	icos_lut[7772] =  9'sd162;
	qsin_lut[7773] = -9'sd127;
	icos_lut[7773] =  9'sd190;
	qsin_lut[7774] = -9'sd88;
	icos_lut[7774] =  9'sd212;
	qsin_lut[7775] = -9'sd45;
	icos_lut[7775] =  9'sd225;
	qsin_lut[7776] =  9'sd0;
	icos_lut[7776] =  9'sd231;
	qsin_lut[7777] =  9'sd45;
	icos_lut[7777] =  9'sd227;
	qsin_lut[7778] =  9'sd88;
	icos_lut[7778] =  9'sd213;
	qsin_lut[7779] =  9'sd128;
	icos_lut[7779] =  9'sd192;
	qsin_lut[7780] =  9'sd163;
	icos_lut[7780] =  9'sd163;
	qsin_lut[7781] =  9'sd192;
	icos_lut[7781] =  9'sd128;
	qsin_lut[7782] =  9'sd213;
	icos_lut[7782] =  9'sd88;
	qsin_lut[7783] =  9'sd227;
	icos_lut[7783] =  9'sd45;
	qsin_lut[7784] =  9'sd231;
	icos_lut[7784] =  9'sd0;
	qsin_lut[7785] =  9'sd227;
	icos_lut[7785] = -9'sd45;
	qsin_lut[7786] =  9'sd213;
	icos_lut[7786] = -9'sd88;
	qsin_lut[7787] =  9'sd192;
	icos_lut[7787] = -9'sd128;
	qsin_lut[7788] =  9'sd163;
	icos_lut[7788] = -9'sd163;
	qsin_lut[7789] =  9'sd128;
	icos_lut[7789] = -9'sd192;
	qsin_lut[7790] =  9'sd88;
	icos_lut[7790] = -9'sd213;
	qsin_lut[7791] =  9'sd45;
	icos_lut[7791] = -9'sd227;
	qsin_lut[7792] =  9'sd0;
	icos_lut[7792] = -9'sd231;
	qsin_lut[7793] = -9'sd45;
	icos_lut[7793] = -9'sd227;
	qsin_lut[7794] = -9'sd88;
	icos_lut[7794] = -9'sd213;
	qsin_lut[7795] = -9'sd128;
	icos_lut[7795] = -9'sd192;
	qsin_lut[7796] = -9'sd163;
	icos_lut[7796] = -9'sd163;
	qsin_lut[7797] = -9'sd192;
	icos_lut[7797] = -9'sd128;
	qsin_lut[7798] = -9'sd213;
	icos_lut[7798] = -9'sd88;
	qsin_lut[7799] = -9'sd227;
	icos_lut[7799] = -9'sd45;
	qsin_lut[7800] = -9'sd231;
	icos_lut[7800] = -9'sd0;
	qsin_lut[7801] = -9'sd227;
	icos_lut[7801] =  9'sd45;
	qsin_lut[7802] = -9'sd213;
	icos_lut[7802] =  9'sd88;
	qsin_lut[7803] = -9'sd192;
	icos_lut[7803] =  9'sd128;
	qsin_lut[7804] = -9'sd163;
	icos_lut[7804] =  9'sd163;
	qsin_lut[7805] = -9'sd128;
	icos_lut[7805] =  9'sd192;
	qsin_lut[7806] = -9'sd88;
	icos_lut[7806] =  9'sd213;
	qsin_lut[7807] = -9'sd45;
	icos_lut[7807] =  9'sd227;
	qsin_lut[7808] =  9'sd0;
	icos_lut[7808] =  9'sd233;
	qsin_lut[7809] =  9'sd45;
	icos_lut[7809] =  9'sd229;
	qsin_lut[7810] =  9'sd89;
	icos_lut[7810] =  9'sd215;
	qsin_lut[7811] =  9'sd129;
	icos_lut[7811] =  9'sd194;
	qsin_lut[7812] =  9'sd165;
	icos_lut[7812] =  9'sd165;
	qsin_lut[7813] =  9'sd194;
	icos_lut[7813] =  9'sd129;
	qsin_lut[7814] =  9'sd215;
	icos_lut[7814] =  9'sd89;
	qsin_lut[7815] =  9'sd229;
	icos_lut[7815] =  9'sd45;
	qsin_lut[7816] =  9'sd233;
	icos_lut[7816] =  9'sd0;
	qsin_lut[7817] =  9'sd229;
	icos_lut[7817] = -9'sd45;
	qsin_lut[7818] =  9'sd215;
	icos_lut[7818] = -9'sd89;
	qsin_lut[7819] =  9'sd194;
	icos_lut[7819] = -9'sd129;
	qsin_lut[7820] =  9'sd165;
	icos_lut[7820] = -9'sd165;
	qsin_lut[7821] =  9'sd129;
	icos_lut[7821] = -9'sd194;
	qsin_lut[7822] =  9'sd89;
	icos_lut[7822] = -9'sd215;
	qsin_lut[7823] =  9'sd45;
	icos_lut[7823] = -9'sd229;
	qsin_lut[7824] =  9'sd0;
	icos_lut[7824] = -9'sd233;
	qsin_lut[7825] = -9'sd45;
	icos_lut[7825] = -9'sd229;
	qsin_lut[7826] = -9'sd89;
	icos_lut[7826] = -9'sd215;
	qsin_lut[7827] = -9'sd129;
	icos_lut[7827] = -9'sd194;
	qsin_lut[7828] = -9'sd165;
	icos_lut[7828] = -9'sd165;
	qsin_lut[7829] = -9'sd194;
	icos_lut[7829] = -9'sd129;
	qsin_lut[7830] = -9'sd215;
	icos_lut[7830] = -9'sd89;
	qsin_lut[7831] = -9'sd229;
	icos_lut[7831] = -9'sd45;
	qsin_lut[7832] = -9'sd233;
	icos_lut[7832] = -9'sd0;
	qsin_lut[7833] = -9'sd229;
	icos_lut[7833] =  9'sd45;
	qsin_lut[7834] = -9'sd215;
	icos_lut[7834] =  9'sd89;
	qsin_lut[7835] = -9'sd194;
	icos_lut[7835] =  9'sd129;
	qsin_lut[7836] = -9'sd165;
	icos_lut[7836] =  9'sd165;
	qsin_lut[7837] = -9'sd129;
	icos_lut[7837] =  9'sd194;
	qsin_lut[7838] = -9'sd89;
	icos_lut[7838] =  9'sd215;
	qsin_lut[7839] = -9'sd45;
	icos_lut[7839] =  9'sd229;
	qsin_lut[7840] =  9'sd0;
	icos_lut[7840] =  9'sd235;
	qsin_lut[7841] =  9'sd46;
	icos_lut[7841] =  9'sd230;
	qsin_lut[7842] =  9'sd90;
	icos_lut[7842] =  9'sd217;
	qsin_lut[7843] =  9'sd131;
	icos_lut[7843] =  9'sd195;
	qsin_lut[7844] =  9'sd166;
	icos_lut[7844] =  9'sd166;
	qsin_lut[7845] =  9'sd195;
	icos_lut[7845] =  9'sd131;
	qsin_lut[7846] =  9'sd217;
	icos_lut[7846] =  9'sd90;
	qsin_lut[7847] =  9'sd230;
	icos_lut[7847] =  9'sd46;
	qsin_lut[7848] =  9'sd235;
	icos_lut[7848] =  9'sd0;
	qsin_lut[7849] =  9'sd230;
	icos_lut[7849] = -9'sd46;
	qsin_lut[7850] =  9'sd217;
	icos_lut[7850] = -9'sd90;
	qsin_lut[7851] =  9'sd195;
	icos_lut[7851] = -9'sd131;
	qsin_lut[7852] =  9'sd166;
	icos_lut[7852] = -9'sd166;
	qsin_lut[7853] =  9'sd131;
	icos_lut[7853] = -9'sd195;
	qsin_lut[7854] =  9'sd90;
	icos_lut[7854] = -9'sd217;
	qsin_lut[7855] =  9'sd46;
	icos_lut[7855] = -9'sd230;
	qsin_lut[7856] =  9'sd0;
	icos_lut[7856] = -9'sd235;
	qsin_lut[7857] = -9'sd46;
	icos_lut[7857] = -9'sd230;
	qsin_lut[7858] = -9'sd90;
	icos_lut[7858] = -9'sd217;
	qsin_lut[7859] = -9'sd131;
	icos_lut[7859] = -9'sd195;
	qsin_lut[7860] = -9'sd166;
	icos_lut[7860] = -9'sd166;
	qsin_lut[7861] = -9'sd195;
	icos_lut[7861] = -9'sd131;
	qsin_lut[7862] = -9'sd217;
	icos_lut[7862] = -9'sd90;
	qsin_lut[7863] = -9'sd230;
	icos_lut[7863] = -9'sd46;
	qsin_lut[7864] = -9'sd235;
	icos_lut[7864] = -9'sd0;
	qsin_lut[7865] = -9'sd230;
	icos_lut[7865] =  9'sd46;
	qsin_lut[7866] = -9'sd217;
	icos_lut[7866] =  9'sd90;
	qsin_lut[7867] = -9'sd195;
	icos_lut[7867] =  9'sd131;
	qsin_lut[7868] = -9'sd166;
	icos_lut[7868] =  9'sd166;
	qsin_lut[7869] = -9'sd131;
	icos_lut[7869] =  9'sd195;
	qsin_lut[7870] = -9'sd90;
	icos_lut[7870] =  9'sd217;
	qsin_lut[7871] = -9'sd46;
	icos_lut[7871] =  9'sd230;
	qsin_lut[7872] =  9'sd0;
	icos_lut[7872] =  9'sd237;
	qsin_lut[7873] =  9'sd46;
	icos_lut[7873] =  9'sd232;
	qsin_lut[7874] =  9'sd91;
	icos_lut[7874] =  9'sd219;
	qsin_lut[7875] =  9'sd132;
	icos_lut[7875] =  9'sd197;
	qsin_lut[7876] =  9'sd168;
	icos_lut[7876] =  9'sd168;
	qsin_lut[7877] =  9'sd197;
	icos_lut[7877] =  9'sd132;
	qsin_lut[7878] =  9'sd219;
	icos_lut[7878] =  9'sd91;
	qsin_lut[7879] =  9'sd232;
	icos_lut[7879] =  9'sd46;
	qsin_lut[7880] =  9'sd237;
	icos_lut[7880] =  9'sd0;
	qsin_lut[7881] =  9'sd232;
	icos_lut[7881] = -9'sd46;
	qsin_lut[7882] =  9'sd219;
	icos_lut[7882] = -9'sd91;
	qsin_lut[7883] =  9'sd197;
	icos_lut[7883] = -9'sd132;
	qsin_lut[7884] =  9'sd168;
	icos_lut[7884] = -9'sd168;
	qsin_lut[7885] =  9'sd132;
	icos_lut[7885] = -9'sd197;
	qsin_lut[7886] =  9'sd91;
	icos_lut[7886] = -9'sd219;
	qsin_lut[7887] =  9'sd46;
	icos_lut[7887] = -9'sd232;
	qsin_lut[7888] =  9'sd0;
	icos_lut[7888] = -9'sd237;
	qsin_lut[7889] = -9'sd46;
	icos_lut[7889] = -9'sd232;
	qsin_lut[7890] = -9'sd91;
	icos_lut[7890] = -9'sd219;
	qsin_lut[7891] = -9'sd132;
	icos_lut[7891] = -9'sd197;
	qsin_lut[7892] = -9'sd168;
	icos_lut[7892] = -9'sd168;
	qsin_lut[7893] = -9'sd197;
	icos_lut[7893] = -9'sd132;
	qsin_lut[7894] = -9'sd219;
	icos_lut[7894] = -9'sd91;
	qsin_lut[7895] = -9'sd232;
	icos_lut[7895] = -9'sd46;
	qsin_lut[7896] = -9'sd237;
	icos_lut[7896] = -9'sd0;
	qsin_lut[7897] = -9'sd232;
	icos_lut[7897] =  9'sd46;
	qsin_lut[7898] = -9'sd219;
	icos_lut[7898] =  9'sd91;
	qsin_lut[7899] = -9'sd197;
	icos_lut[7899] =  9'sd132;
	qsin_lut[7900] = -9'sd168;
	icos_lut[7900] =  9'sd168;
	qsin_lut[7901] = -9'sd132;
	icos_lut[7901] =  9'sd197;
	qsin_lut[7902] = -9'sd91;
	icos_lut[7902] =  9'sd219;
	qsin_lut[7903] = -9'sd46;
	icos_lut[7903] =  9'sd232;
	qsin_lut[7904] =  9'sd0;
	icos_lut[7904] =  9'sd239;
	qsin_lut[7905] =  9'sd47;
	icos_lut[7905] =  9'sd234;
	qsin_lut[7906] =  9'sd91;
	icos_lut[7906] =  9'sd221;
	qsin_lut[7907] =  9'sd133;
	icos_lut[7907] =  9'sd199;
	qsin_lut[7908] =  9'sd169;
	icos_lut[7908] =  9'sd169;
	qsin_lut[7909] =  9'sd199;
	icos_lut[7909] =  9'sd133;
	qsin_lut[7910] =  9'sd221;
	icos_lut[7910] =  9'sd91;
	qsin_lut[7911] =  9'sd234;
	icos_lut[7911] =  9'sd47;
	qsin_lut[7912] =  9'sd239;
	icos_lut[7912] =  9'sd0;
	qsin_lut[7913] =  9'sd234;
	icos_lut[7913] = -9'sd47;
	qsin_lut[7914] =  9'sd221;
	icos_lut[7914] = -9'sd91;
	qsin_lut[7915] =  9'sd199;
	icos_lut[7915] = -9'sd133;
	qsin_lut[7916] =  9'sd169;
	icos_lut[7916] = -9'sd169;
	qsin_lut[7917] =  9'sd133;
	icos_lut[7917] = -9'sd199;
	qsin_lut[7918] =  9'sd91;
	icos_lut[7918] = -9'sd221;
	qsin_lut[7919] =  9'sd47;
	icos_lut[7919] = -9'sd234;
	qsin_lut[7920] =  9'sd0;
	icos_lut[7920] = -9'sd239;
	qsin_lut[7921] = -9'sd47;
	icos_lut[7921] = -9'sd234;
	qsin_lut[7922] = -9'sd91;
	icos_lut[7922] = -9'sd221;
	qsin_lut[7923] = -9'sd133;
	icos_lut[7923] = -9'sd199;
	qsin_lut[7924] = -9'sd169;
	icos_lut[7924] = -9'sd169;
	qsin_lut[7925] = -9'sd199;
	icos_lut[7925] = -9'sd133;
	qsin_lut[7926] = -9'sd221;
	icos_lut[7926] = -9'sd91;
	qsin_lut[7927] = -9'sd234;
	icos_lut[7927] = -9'sd47;
	qsin_lut[7928] = -9'sd239;
	icos_lut[7928] = -9'sd0;
	qsin_lut[7929] = -9'sd234;
	icos_lut[7929] =  9'sd47;
	qsin_lut[7930] = -9'sd221;
	icos_lut[7930] =  9'sd91;
	qsin_lut[7931] = -9'sd199;
	icos_lut[7931] =  9'sd133;
	qsin_lut[7932] = -9'sd169;
	icos_lut[7932] =  9'sd169;
	qsin_lut[7933] = -9'sd133;
	icos_lut[7933] =  9'sd199;
	qsin_lut[7934] = -9'sd91;
	icos_lut[7934] =  9'sd221;
	qsin_lut[7935] = -9'sd47;
	icos_lut[7935] =  9'sd234;
	qsin_lut[7936] =  9'sd0;
	icos_lut[7936] =  9'sd241;
	qsin_lut[7937] =  9'sd47;
	icos_lut[7937] =  9'sd236;
	qsin_lut[7938] =  9'sd92;
	icos_lut[7938] =  9'sd223;
	qsin_lut[7939] =  9'sd134;
	icos_lut[7939] =  9'sd200;
	qsin_lut[7940] =  9'sd170;
	icos_lut[7940] =  9'sd170;
	qsin_lut[7941] =  9'sd200;
	icos_lut[7941] =  9'sd134;
	qsin_lut[7942] =  9'sd223;
	icos_lut[7942] =  9'sd92;
	qsin_lut[7943] =  9'sd236;
	icos_lut[7943] =  9'sd47;
	qsin_lut[7944] =  9'sd241;
	icos_lut[7944] =  9'sd0;
	qsin_lut[7945] =  9'sd236;
	icos_lut[7945] = -9'sd47;
	qsin_lut[7946] =  9'sd223;
	icos_lut[7946] = -9'sd92;
	qsin_lut[7947] =  9'sd200;
	icos_lut[7947] = -9'sd134;
	qsin_lut[7948] =  9'sd170;
	icos_lut[7948] = -9'sd170;
	qsin_lut[7949] =  9'sd134;
	icos_lut[7949] = -9'sd200;
	qsin_lut[7950] =  9'sd92;
	icos_lut[7950] = -9'sd223;
	qsin_lut[7951] =  9'sd47;
	icos_lut[7951] = -9'sd236;
	qsin_lut[7952] =  9'sd0;
	icos_lut[7952] = -9'sd241;
	qsin_lut[7953] = -9'sd47;
	icos_lut[7953] = -9'sd236;
	qsin_lut[7954] = -9'sd92;
	icos_lut[7954] = -9'sd223;
	qsin_lut[7955] = -9'sd134;
	icos_lut[7955] = -9'sd200;
	qsin_lut[7956] = -9'sd170;
	icos_lut[7956] = -9'sd170;
	qsin_lut[7957] = -9'sd200;
	icos_lut[7957] = -9'sd134;
	qsin_lut[7958] = -9'sd223;
	icos_lut[7958] = -9'sd92;
	qsin_lut[7959] = -9'sd236;
	icos_lut[7959] = -9'sd47;
	qsin_lut[7960] = -9'sd241;
	icos_lut[7960] = -9'sd0;
	qsin_lut[7961] = -9'sd236;
	icos_lut[7961] =  9'sd47;
	qsin_lut[7962] = -9'sd223;
	icos_lut[7962] =  9'sd92;
	qsin_lut[7963] = -9'sd200;
	icos_lut[7963] =  9'sd134;
	qsin_lut[7964] = -9'sd170;
	icos_lut[7964] =  9'sd170;
	qsin_lut[7965] = -9'sd134;
	icos_lut[7965] =  9'sd200;
	qsin_lut[7966] = -9'sd92;
	icos_lut[7966] =  9'sd223;
	qsin_lut[7967] = -9'sd47;
	icos_lut[7967] =  9'sd236;
	qsin_lut[7968] =  9'sd0;
	icos_lut[7968] =  9'sd243;
	qsin_lut[7969] =  9'sd47;
	icos_lut[7969] =  9'sd238;
	qsin_lut[7970] =  9'sd93;
	icos_lut[7970] =  9'sd225;
	qsin_lut[7971] =  9'sd135;
	icos_lut[7971] =  9'sd202;
	qsin_lut[7972] =  9'sd172;
	icos_lut[7972] =  9'sd172;
	qsin_lut[7973] =  9'sd202;
	icos_lut[7973] =  9'sd135;
	qsin_lut[7974] =  9'sd225;
	icos_lut[7974] =  9'sd93;
	qsin_lut[7975] =  9'sd238;
	icos_lut[7975] =  9'sd47;
	qsin_lut[7976] =  9'sd243;
	icos_lut[7976] =  9'sd0;
	qsin_lut[7977] =  9'sd238;
	icos_lut[7977] = -9'sd47;
	qsin_lut[7978] =  9'sd225;
	icos_lut[7978] = -9'sd93;
	qsin_lut[7979] =  9'sd202;
	icos_lut[7979] = -9'sd135;
	qsin_lut[7980] =  9'sd172;
	icos_lut[7980] = -9'sd172;
	qsin_lut[7981] =  9'sd135;
	icos_lut[7981] = -9'sd202;
	qsin_lut[7982] =  9'sd93;
	icos_lut[7982] = -9'sd225;
	qsin_lut[7983] =  9'sd47;
	icos_lut[7983] = -9'sd238;
	qsin_lut[7984] =  9'sd0;
	icos_lut[7984] = -9'sd243;
	qsin_lut[7985] = -9'sd47;
	icos_lut[7985] = -9'sd238;
	qsin_lut[7986] = -9'sd93;
	icos_lut[7986] = -9'sd225;
	qsin_lut[7987] = -9'sd135;
	icos_lut[7987] = -9'sd202;
	qsin_lut[7988] = -9'sd172;
	icos_lut[7988] = -9'sd172;
	qsin_lut[7989] = -9'sd202;
	icos_lut[7989] = -9'sd135;
	qsin_lut[7990] = -9'sd225;
	icos_lut[7990] = -9'sd93;
	qsin_lut[7991] = -9'sd238;
	icos_lut[7991] = -9'sd47;
	qsin_lut[7992] = -9'sd243;
	icos_lut[7992] = -9'sd0;
	qsin_lut[7993] = -9'sd238;
	icos_lut[7993] =  9'sd47;
	qsin_lut[7994] = -9'sd225;
	icos_lut[7994] =  9'sd93;
	qsin_lut[7995] = -9'sd202;
	icos_lut[7995] =  9'sd135;
	qsin_lut[7996] = -9'sd172;
	icos_lut[7996] =  9'sd172;
	qsin_lut[7997] = -9'sd135;
	icos_lut[7997] =  9'sd202;
	qsin_lut[7998] = -9'sd93;
	icos_lut[7998] =  9'sd225;
	qsin_lut[7999] = -9'sd47;
	icos_lut[7999] =  9'sd238;
	qsin_lut[8000] =  9'sd0;
	icos_lut[8000] =  9'sd245;
	qsin_lut[8001] =  9'sd48;
	icos_lut[8001] =  9'sd240;
	qsin_lut[8002] =  9'sd94;
	icos_lut[8002] =  9'sd226;
	qsin_lut[8003] =  9'sd136;
	icos_lut[8003] =  9'sd204;
	qsin_lut[8004] =  9'sd173;
	icos_lut[8004] =  9'sd173;
	qsin_lut[8005] =  9'sd204;
	icos_lut[8005] =  9'sd136;
	qsin_lut[8006] =  9'sd226;
	icos_lut[8006] =  9'sd94;
	qsin_lut[8007] =  9'sd240;
	icos_lut[8007] =  9'sd48;
	qsin_lut[8008] =  9'sd245;
	icos_lut[8008] =  9'sd0;
	qsin_lut[8009] =  9'sd240;
	icos_lut[8009] = -9'sd48;
	qsin_lut[8010] =  9'sd226;
	icos_lut[8010] = -9'sd94;
	qsin_lut[8011] =  9'sd204;
	icos_lut[8011] = -9'sd136;
	qsin_lut[8012] =  9'sd173;
	icos_lut[8012] = -9'sd173;
	qsin_lut[8013] =  9'sd136;
	icos_lut[8013] = -9'sd204;
	qsin_lut[8014] =  9'sd94;
	icos_lut[8014] = -9'sd226;
	qsin_lut[8015] =  9'sd48;
	icos_lut[8015] = -9'sd240;
	qsin_lut[8016] =  9'sd0;
	icos_lut[8016] = -9'sd245;
	qsin_lut[8017] = -9'sd48;
	icos_lut[8017] = -9'sd240;
	qsin_lut[8018] = -9'sd94;
	icos_lut[8018] = -9'sd226;
	qsin_lut[8019] = -9'sd136;
	icos_lut[8019] = -9'sd204;
	qsin_lut[8020] = -9'sd173;
	icos_lut[8020] = -9'sd173;
	qsin_lut[8021] = -9'sd204;
	icos_lut[8021] = -9'sd136;
	qsin_lut[8022] = -9'sd226;
	icos_lut[8022] = -9'sd94;
	qsin_lut[8023] = -9'sd240;
	icos_lut[8023] = -9'sd48;
	qsin_lut[8024] = -9'sd245;
	icos_lut[8024] = -9'sd0;
	qsin_lut[8025] = -9'sd240;
	icos_lut[8025] =  9'sd48;
	qsin_lut[8026] = -9'sd226;
	icos_lut[8026] =  9'sd94;
	qsin_lut[8027] = -9'sd204;
	icos_lut[8027] =  9'sd136;
	qsin_lut[8028] = -9'sd173;
	icos_lut[8028] =  9'sd173;
	qsin_lut[8029] = -9'sd136;
	icos_lut[8029] =  9'sd204;
	qsin_lut[8030] = -9'sd94;
	icos_lut[8030] =  9'sd226;
	qsin_lut[8031] = -9'sd48;
	icos_lut[8031] =  9'sd240;
	qsin_lut[8032] =  9'sd0;
	icos_lut[8032] =  9'sd247;
	qsin_lut[8033] =  9'sd48;
	icos_lut[8033] =  9'sd242;
	qsin_lut[8034] =  9'sd95;
	icos_lut[8034] =  9'sd228;
	qsin_lut[8035] =  9'sd137;
	icos_lut[8035] =  9'sd205;
	qsin_lut[8036] =  9'sd175;
	icos_lut[8036] =  9'sd175;
	qsin_lut[8037] =  9'sd205;
	icos_lut[8037] =  9'sd137;
	qsin_lut[8038] =  9'sd228;
	icos_lut[8038] =  9'sd95;
	qsin_lut[8039] =  9'sd242;
	icos_lut[8039] =  9'sd48;
	qsin_lut[8040] =  9'sd247;
	icos_lut[8040] =  9'sd0;
	qsin_lut[8041] =  9'sd242;
	icos_lut[8041] = -9'sd48;
	qsin_lut[8042] =  9'sd228;
	icos_lut[8042] = -9'sd95;
	qsin_lut[8043] =  9'sd205;
	icos_lut[8043] = -9'sd137;
	qsin_lut[8044] =  9'sd175;
	icos_lut[8044] = -9'sd175;
	qsin_lut[8045] =  9'sd137;
	icos_lut[8045] = -9'sd205;
	qsin_lut[8046] =  9'sd95;
	icos_lut[8046] = -9'sd228;
	qsin_lut[8047] =  9'sd48;
	icos_lut[8047] = -9'sd242;
	qsin_lut[8048] =  9'sd0;
	icos_lut[8048] = -9'sd247;
	qsin_lut[8049] = -9'sd48;
	icos_lut[8049] = -9'sd242;
	qsin_lut[8050] = -9'sd95;
	icos_lut[8050] = -9'sd228;
	qsin_lut[8051] = -9'sd137;
	icos_lut[8051] = -9'sd205;
	qsin_lut[8052] = -9'sd175;
	icos_lut[8052] = -9'sd175;
	qsin_lut[8053] = -9'sd205;
	icos_lut[8053] = -9'sd137;
	qsin_lut[8054] = -9'sd228;
	icos_lut[8054] = -9'sd95;
	qsin_lut[8055] = -9'sd242;
	icos_lut[8055] = -9'sd48;
	qsin_lut[8056] = -9'sd247;
	icos_lut[8056] = -9'sd0;
	qsin_lut[8057] = -9'sd242;
	icos_lut[8057] =  9'sd48;
	qsin_lut[8058] = -9'sd228;
	icos_lut[8058] =  9'sd95;
	qsin_lut[8059] = -9'sd205;
	icos_lut[8059] =  9'sd137;
	qsin_lut[8060] = -9'sd175;
	icos_lut[8060] =  9'sd175;
	qsin_lut[8061] = -9'sd137;
	icos_lut[8061] =  9'sd205;
	qsin_lut[8062] = -9'sd95;
	icos_lut[8062] =  9'sd228;
	qsin_lut[8063] = -9'sd48;
	icos_lut[8063] =  9'sd242;
	qsin_lut[8064] =  9'sd0;
	icos_lut[8064] =  9'sd249;
	qsin_lut[8065] =  9'sd49;
	icos_lut[8065] =  9'sd244;
	qsin_lut[8066] =  9'sd95;
	icos_lut[8066] =  9'sd230;
	qsin_lut[8067] =  9'sd138;
	icos_lut[8067] =  9'sd207;
	qsin_lut[8068] =  9'sd176;
	icos_lut[8068] =  9'sd176;
	qsin_lut[8069] =  9'sd207;
	icos_lut[8069] =  9'sd138;
	qsin_lut[8070] =  9'sd230;
	icos_lut[8070] =  9'sd95;
	qsin_lut[8071] =  9'sd244;
	icos_lut[8071] =  9'sd49;
	qsin_lut[8072] =  9'sd249;
	icos_lut[8072] =  9'sd0;
	qsin_lut[8073] =  9'sd244;
	icos_lut[8073] = -9'sd49;
	qsin_lut[8074] =  9'sd230;
	icos_lut[8074] = -9'sd95;
	qsin_lut[8075] =  9'sd207;
	icos_lut[8075] = -9'sd138;
	qsin_lut[8076] =  9'sd176;
	icos_lut[8076] = -9'sd176;
	qsin_lut[8077] =  9'sd138;
	icos_lut[8077] = -9'sd207;
	qsin_lut[8078] =  9'sd95;
	icos_lut[8078] = -9'sd230;
	qsin_lut[8079] =  9'sd49;
	icos_lut[8079] = -9'sd244;
	qsin_lut[8080] =  9'sd0;
	icos_lut[8080] = -9'sd249;
	qsin_lut[8081] = -9'sd49;
	icos_lut[8081] = -9'sd244;
	qsin_lut[8082] = -9'sd95;
	icos_lut[8082] = -9'sd230;
	qsin_lut[8083] = -9'sd138;
	icos_lut[8083] = -9'sd207;
	qsin_lut[8084] = -9'sd176;
	icos_lut[8084] = -9'sd176;
	qsin_lut[8085] = -9'sd207;
	icos_lut[8085] = -9'sd138;
	qsin_lut[8086] = -9'sd230;
	icos_lut[8086] = -9'sd95;
	qsin_lut[8087] = -9'sd244;
	icos_lut[8087] = -9'sd49;
	qsin_lut[8088] = -9'sd249;
	icos_lut[8088] = -9'sd0;
	qsin_lut[8089] = -9'sd244;
	icos_lut[8089] =  9'sd49;
	qsin_lut[8090] = -9'sd230;
	icos_lut[8090] =  9'sd95;
	qsin_lut[8091] = -9'sd207;
	icos_lut[8091] =  9'sd138;
	qsin_lut[8092] = -9'sd176;
	icos_lut[8092] =  9'sd176;
	qsin_lut[8093] = -9'sd138;
	icos_lut[8093] =  9'sd207;
	qsin_lut[8094] = -9'sd95;
	icos_lut[8094] =  9'sd230;
	qsin_lut[8095] = -9'sd49;
	icos_lut[8095] =  9'sd244;
	qsin_lut[8096] =  9'sd0;
	icos_lut[8096] =  9'sd251;
	qsin_lut[8097] =  9'sd49;
	icos_lut[8097] =  9'sd246;
	qsin_lut[8098] =  9'sd96;
	icos_lut[8098] =  9'sd232;
	qsin_lut[8099] =  9'sd139;
	icos_lut[8099] =  9'sd209;
	qsin_lut[8100] =  9'sd177;
	icos_lut[8100] =  9'sd177;
	qsin_lut[8101] =  9'sd209;
	icos_lut[8101] =  9'sd139;
	qsin_lut[8102] =  9'sd232;
	icos_lut[8102] =  9'sd96;
	qsin_lut[8103] =  9'sd246;
	icos_lut[8103] =  9'sd49;
	qsin_lut[8104] =  9'sd251;
	icos_lut[8104] =  9'sd0;
	qsin_lut[8105] =  9'sd246;
	icos_lut[8105] = -9'sd49;
	qsin_lut[8106] =  9'sd232;
	icos_lut[8106] = -9'sd96;
	qsin_lut[8107] =  9'sd209;
	icos_lut[8107] = -9'sd139;
	qsin_lut[8108] =  9'sd177;
	icos_lut[8108] = -9'sd177;
	qsin_lut[8109] =  9'sd139;
	icos_lut[8109] = -9'sd209;
	qsin_lut[8110] =  9'sd96;
	icos_lut[8110] = -9'sd232;
	qsin_lut[8111] =  9'sd49;
	icos_lut[8111] = -9'sd246;
	qsin_lut[8112] =  9'sd0;
	icos_lut[8112] = -9'sd251;
	qsin_lut[8113] = -9'sd49;
	icos_lut[8113] = -9'sd246;
	qsin_lut[8114] = -9'sd96;
	icos_lut[8114] = -9'sd232;
	qsin_lut[8115] = -9'sd139;
	icos_lut[8115] = -9'sd209;
	qsin_lut[8116] = -9'sd177;
	icos_lut[8116] = -9'sd177;
	qsin_lut[8117] = -9'sd209;
	icos_lut[8117] = -9'sd139;
	qsin_lut[8118] = -9'sd232;
	icos_lut[8118] = -9'sd96;
	qsin_lut[8119] = -9'sd246;
	icos_lut[8119] = -9'sd49;
	qsin_lut[8120] = -9'sd251;
	icos_lut[8120] = -9'sd0;
	qsin_lut[8121] = -9'sd246;
	icos_lut[8121] =  9'sd49;
	qsin_lut[8122] = -9'sd232;
	icos_lut[8122] =  9'sd96;
	qsin_lut[8123] = -9'sd209;
	icos_lut[8123] =  9'sd139;
	qsin_lut[8124] = -9'sd177;
	icos_lut[8124] =  9'sd177;
	qsin_lut[8125] = -9'sd139;
	icos_lut[8125] =  9'sd209;
	qsin_lut[8126] = -9'sd96;
	icos_lut[8126] =  9'sd232;
	qsin_lut[8127] = -9'sd49;
	icos_lut[8127] =  9'sd246;
	qsin_lut[8128] =  9'sd0;
	icos_lut[8128] =  9'sd253;
	qsin_lut[8129] =  9'sd49;
	icos_lut[8129] =  9'sd248;
	qsin_lut[8130] =  9'sd97;
	icos_lut[8130] =  9'sd234;
	qsin_lut[8131] =  9'sd141;
	icos_lut[8131] =  9'sd210;
	qsin_lut[8132] =  9'sd179;
	icos_lut[8132] =  9'sd179;
	qsin_lut[8133] =  9'sd210;
	icos_lut[8133] =  9'sd141;
	qsin_lut[8134] =  9'sd234;
	icos_lut[8134] =  9'sd97;
	qsin_lut[8135] =  9'sd248;
	icos_lut[8135] =  9'sd49;
	qsin_lut[8136] =  9'sd253;
	icos_lut[8136] =  9'sd0;
	qsin_lut[8137] =  9'sd248;
	icos_lut[8137] = -9'sd49;
	qsin_lut[8138] =  9'sd234;
	icos_lut[8138] = -9'sd97;
	qsin_lut[8139] =  9'sd210;
	icos_lut[8139] = -9'sd141;
	qsin_lut[8140] =  9'sd179;
	icos_lut[8140] = -9'sd179;
	qsin_lut[8141] =  9'sd141;
	icos_lut[8141] = -9'sd210;
	qsin_lut[8142] =  9'sd97;
	icos_lut[8142] = -9'sd234;
	qsin_lut[8143] =  9'sd49;
	icos_lut[8143] = -9'sd248;
	qsin_lut[8144] =  9'sd0;
	icos_lut[8144] = -9'sd253;
	qsin_lut[8145] = -9'sd49;
	icos_lut[8145] = -9'sd248;
	qsin_lut[8146] = -9'sd97;
	icos_lut[8146] = -9'sd234;
	qsin_lut[8147] = -9'sd141;
	icos_lut[8147] = -9'sd210;
	qsin_lut[8148] = -9'sd179;
	icos_lut[8148] = -9'sd179;
	qsin_lut[8149] = -9'sd210;
	icos_lut[8149] = -9'sd141;
	qsin_lut[8150] = -9'sd234;
	icos_lut[8150] = -9'sd97;
	qsin_lut[8151] = -9'sd248;
	icos_lut[8151] = -9'sd49;
	qsin_lut[8152] = -9'sd253;
	icos_lut[8152] = -9'sd0;
	qsin_lut[8153] = -9'sd248;
	icos_lut[8153] =  9'sd49;
	qsin_lut[8154] = -9'sd234;
	icos_lut[8154] =  9'sd97;
	qsin_lut[8155] = -9'sd210;
	icos_lut[8155] =  9'sd141;
	qsin_lut[8156] = -9'sd179;
	icos_lut[8156] =  9'sd179;
	qsin_lut[8157] = -9'sd141;
	icos_lut[8157] =  9'sd210;
	qsin_lut[8158] = -9'sd97;
	icos_lut[8158] =  9'sd234;
	qsin_lut[8159] = -9'sd49;
	icos_lut[8159] =  9'sd248;
	qsin_lut[8160] =  9'sd0;
	icos_lut[8160] =  9'sd255;
	qsin_lut[8161] =  9'sd50;
	icos_lut[8161] =  9'sd250;
	qsin_lut[8162] =  9'sd98;
	icos_lut[8162] =  9'sd236;
	qsin_lut[8163] =  9'sd142;
	icos_lut[8163] =  9'sd212;
	qsin_lut[8164] =  9'sd180;
	icos_lut[8164] =  9'sd180;
	qsin_lut[8165] =  9'sd212;
	icos_lut[8165] =  9'sd142;
	qsin_lut[8166] =  9'sd236;
	icos_lut[8166] =  9'sd98;
	qsin_lut[8167] =  9'sd250;
	icos_lut[8167] =  9'sd50;
	qsin_lut[8168] =  9'sd255;
	icos_lut[8168] =  9'sd0;
	qsin_lut[8169] =  9'sd250;
	icos_lut[8169] = -9'sd50;
	qsin_lut[8170] =  9'sd236;
	icos_lut[8170] = -9'sd98;
	qsin_lut[8171] =  9'sd212;
	icos_lut[8171] = -9'sd142;
	qsin_lut[8172] =  9'sd180;
	icos_lut[8172] = -9'sd180;
	qsin_lut[8173] =  9'sd142;
	icos_lut[8173] = -9'sd212;
	qsin_lut[8174] =  9'sd98;
	icos_lut[8174] = -9'sd236;
	qsin_lut[8175] =  9'sd50;
	icos_lut[8175] = -9'sd250;
	qsin_lut[8176] =  9'sd0;
	icos_lut[8176] = -9'sd255;
	qsin_lut[8177] = -9'sd50;
	icos_lut[8177] = -9'sd250;
	qsin_lut[8178] = -9'sd98;
	icos_lut[8178] = -9'sd236;
	qsin_lut[8179] = -9'sd142;
	icos_lut[8179] = -9'sd212;
	qsin_lut[8180] = -9'sd180;
	icos_lut[8180] = -9'sd180;
	qsin_lut[8181] = -9'sd212;
	icos_lut[8181] = -9'sd142;
	qsin_lut[8182] = -9'sd236;
	icos_lut[8182] = -9'sd98;
	qsin_lut[8183] = -9'sd250;
	icos_lut[8183] = -9'sd50;
	qsin_lut[8184] = -9'sd255;
	icos_lut[8184] = -9'sd0;
	qsin_lut[8185] = -9'sd250;
	icos_lut[8185] =  9'sd50;
	qsin_lut[8186] = -9'sd236;
	icos_lut[8186] =  9'sd98;
	qsin_lut[8187] = -9'sd212;
	icos_lut[8187] =  9'sd142;
	qsin_lut[8188] = -9'sd180;
	icos_lut[8188] =  9'sd180;
	qsin_lut[8189] = -9'sd142;
	icos_lut[8189] =  9'sd212;
	qsin_lut[8190] = -9'sd98;
	icos_lut[8190] =  9'sd236;
	qsin_lut[8191] = -9'sd50;
	icos_lut[8191] =  9'sd250;
end
endmodule
