module sincos (
	icos,  //out
	qsin,  //out
	t,	   //in
	i,
	q
);

output [8:0] icos;
output [8:0] qsin;

input [4:0] t;
input [3:0] i;
input [3:0] q;

reg signed [8:0] icos_lut [0:511];
reg signed [8:0] qsin_lut [0:511];

reg [8:0] icos_addr=0;
reg [8:0] qsin_addr=0;
wire [8:0] icos=icos_lut[icos_addr];
wire [8:0] qsin=qsin_lut[qsin_addr];

// address [8:5] is the multiplier, 0:-1, (7,8)=~0, 15=1
// address [4:0] is t

// generated with iq_lut.pl
initial begin
	qsin_lut[000] =  9'sd0;
	icos_lut[000] = -9'sd255;
	qsin_lut[001] = -9'sd50;
	icos_lut[001] = -9'sd250;
	qsin_lut[002] = -9'sd98;
	icos_lut[002] = -9'sd236;
	qsin_lut[003] = -9'sd142;
	icos_lut[003] = -9'sd212;
	qsin_lut[004] = -9'sd180;
	icos_lut[004] = -9'sd180;
	qsin_lut[005] = -9'sd212;
	icos_lut[005] = -9'sd142;
	qsin_lut[006] = -9'sd236;
	icos_lut[006] = -9'sd98;
	qsin_lut[007] = -9'sd250;
	icos_lut[007] = -9'sd50;
	qsin_lut[008] = -9'sd255;
	icos_lut[008] = -9'sd0;
	qsin_lut[009] = -9'sd250;
	icos_lut[009] =  9'sd50;
	qsin_lut[010] = -9'sd236;
	icos_lut[010] =  9'sd98;
	qsin_lut[011] = -9'sd212;
	icos_lut[011] =  9'sd142;
	qsin_lut[012] = -9'sd180;
	icos_lut[012] =  9'sd180;
	qsin_lut[013] = -9'sd142;
	icos_lut[013] =  9'sd212;
	qsin_lut[014] = -9'sd98;
	icos_lut[014] =  9'sd236;
	qsin_lut[015] = -9'sd50;
	icos_lut[015] =  9'sd250;
	qsin_lut[016] = -9'sd0;
	icos_lut[016] =  9'sd255;
	qsin_lut[017] =  9'sd50;
	icos_lut[017] =  9'sd250;
	qsin_lut[018] =  9'sd98;
	icos_lut[018] =  9'sd236;
	qsin_lut[019] =  9'sd142;
	icos_lut[019] =  9'sd212;
	qsin_lut[020] =  9'sd180;
	icos_lut[020] =  9'sd180;
	qsin_lut[021] =  9'sd212;
	icos_lut[021] =  9'sd142;
	qsin_lut[022] =  9'sd236;
	icos_lut[022] =  9'sd98;
	qsin_lut[023] =  9'sd250;
	icos_lut[023] =  9'sd50;
	qsin_lut[024] =  9'sd255;
	icos_lut[024] =  9'sd0;
	qsin_lut[025] =  9'sd250;
	icos_lut[025] = -9'sd50;
	qsin_lut[026] =  9'sd236;
	icos_lut[026] = -9'sd98;
	qsin_lut[027] =  9'sd212;
	icos_lut[027] = -9'sd142;
	qsin_lut[028] =  9'sd180;
	icos_lut[028] = -9'sd180;
	qsin_lut[029] =  9'sd142;
	icos_lut[029] = -9'sd212;
	qsin_lut[030] =  9'sd98;
	icos_lut[030] = -9'sd236;
	qsin_lut[031] =  9'sd50;
	icos_lut[031] = -9'sd250;
	qsin_lut[032] =  9'sd0;
	icos_lut[032] = -9'sd221;
	qsin_lut[033] = -9'sd43;
	icos_lut[033] = -9'sd217;
	qsin_lut[034] = -9'sd85;
	icos_lut[034] = -9'sd204;
	qsin_lut[035] = -9'sd123;
	icos_lut[035] = -9'sd184;
	qsin_lut[036] = -9'sd156;
	icos_lut[036] = -9'sd156;
	qsin_lut[037] = -9'sd184;
	icos_lut[037] = -9'sd123;
	qsin_lut[038] = -9'sd204;
	icos_lut[038] = -9'sd85;
	qsin_lut[039] = -9'sd217;
	icos_lut[039] = -9'sd43;
	qsin_lut[040] = -9'sd221;
	icos_lut[040] = -9'sd0;
	qsin_lut[041] = -9'sd217;
	icos_lut[041] =  9'sd43;
	qsin_lut[042] = -9'sd204;
	icos_lut[042] =  9'sd85;
	qsin_lut[043] = -9'sd184;
	icos_lut[043] =  9'sd123;
	qsin_lut[044] = -9'sd156;
	icos_lut[044] =  9'sd156;
	qsin_lut[045] = -9'sd123;
	icos_lut[045] =  9'sd184;
	qsin_lut[046] = -9'sd85;
	icos_lut[046] =  9'sd204;
	qsin_lut[047] = -9'sd43;
	icos_lut[047] =  9'sd217;
	qsin_lut[048] = -9'sd0;
	icos_lut[048] =  9'sd221;
	qsin_lut[049] =  9'sd43;
	icos_lut[049] =  9'sd217;
	qsin_lut[050] =  9'sd85;
	icos_lut[050] =  9'sd204;
	qsin_lut[051] =  9'sd123;
	icos_lut[051] =  9'sd184;
	qsin_lut[052] =  9'sd156;
	icos_lut[052] =  9'sd156;
	qsin_lut[053] =  9'sd184;
	icos_lut[053] =  9'sd123;
	qsin_lut[054] =  9'sd204;
	icos_lut[054] =  9'sd85;
	qsin_lut[055] =  9'sd217;
	icos_lut[055] =  9'sd43;
	qsin_lut[056] =  9'sd221;
	icos_lut[056] =  9'sd0;
	qsin_lut[057] =  9'sd217;
	icos_lut[057] = -9'sd43;
	qsin_lut[058] =  9'sd204;
	icos_lut[058] = -9'sd85;
	qsin_lut[059] =  9'sd184;
	icos_lut[059] = -9'sd123;
	qsin_lut[060] =  9'sd156;
	icos_lut[060] = -9'sd156;
	qsin_lut[061] =  9'sd123;
	icos_lut[061] = -9'sd184;
	qsin_lut[062] =  9'sd85;
	icos_lut[062] = -9'sd204;
	qsin_lut[063] =  9'sd43;
	icos_lut[063] = -9'sd217;
	qsin_lut[064] =  9'sd0;
	icos_lut[064] = -9'sd187;
	qsin_lut[065] = -9'sd36;
	icos_lut[065] = -9'sd183;
	qsin_lut[066] = -9'sd72;
	icos_lut[066] = -9'sd173;
	qsin_lut[067] = -9'sd104;
	icos_lut[067] = -9'sd155;
	qsin_lut[068] = -9'sd132;
	icos_lut[068] = -9'sd132;
	qsin_lut[069] = -9'sd155;
	icos_lut[069] = -9'sd104;
	qsin_lut[070] = -9'sd173;
	icos_lut[070] = -9'sd72;
	qsin_lut[071] = -9'sd183;
	icos_lut[071] = -9'sd36;
	qsin_lut[072] = -9'sd187;
	icos_lut[072] = -9'sd0;
	qsin_lut[073] = -9'sd183;
	icos_lut[073] =  9'sd36;
	qsin_lut[074] = -9'sd173;
	icos_lut[074] =  9'sd72;
	qsin_lut[075] = -9'sd155;
	icos_lut[075] =  9'sd104;
	qsin_lut[076] = -9'sd132;
	icos_lut[076] =  9'sd132;
	qsin_lut[077] = -9'sd104;
	icos_lut[077] =  9'sd155;
	qsin_lut[078] = -9'sd72;
	icos_lut[078] =  9'sd173;
	qsin_lut[079] = -9'sd36;
	icos_lut[079] =  9'sd183;
	qsin_lut[080] = -9'sd0;
	icos_lut[080] =  9'sd187;
	qsin_lut[081] =  9'sd36;
	icos_lut[081] =  9'sd183;
	qsin_lut[082] =  9'sd72;
	icos_lut[082] =  9'sd173;
	qsin_lut[083] =  9'sd104;
	icos_lut[083] =  9'sd155;
	qsin_lut[084] =  9'sd132;
	icos_lut[084] =  9'sd132;
	qsin_lut[085] =  9'sd155;
	icos_lut[085] =  9'sd104;
	qsin_lut[086] =  9'sd173;
	icos_lut[086] =  9'sd72;
	qsin_lut[087] =  9'sd183;
	icos_lut[087] =  9'sd36;
	qsin_lut[088] =  9'sd187;
	icos_lut[088] =  9'sd0;
	qsin_lut[089] =  9'sd183;
	icos_lut[089] = -9'sd36;
	qsin_lut[090] =  9'sd173;
	icos_lut[090] = -9'sd72;
	qsin_lut[091] =  9'sd155;
	icos_lut[091] = -9'sd104;
	qsin_lut[092] =  9'sd132;
	icos_lut[092] = -9'sd132;
	qsin_lut[093] =  9'sd104;
	icos_lut[093] = -9'sd155;
	qsin_lut[094] =  9'sd72;
	icos_lut[094] = -9'sd173;
	qsin_lut[095] =  9'sd36;
	icos_lut[095] = -9'sd183;
	qsin_lut[096] =  9'sd0;
	icos_lut[096] = -9'sd153;
	qsin_lut[097] = -9'sd30;
	icos_lut[097] = -9'sd150;
	qsin_lut[098] = -9'sd59;
	icos_lut[098] = -9'sd141;
	qsin_lut[099] = -9'sd85;
	icos_lut[099] = -9'sd127;
	qsin_lut[100] = -9'sd108;
	icos_lut[100] = -9'sd108;
	qsin_lut[101] = -9'sd127;
	icos_lut[101] = -9'sd85;
	qsin_lut[102] = -9'sd141;
	icos_lut[102] = -9'sd59;
	qsin_lut[103] = -9'sd150;
	icos_lut[103] = -9'sd30;
	qsin_lut[104] = -9'sd153;
	icos_lut[104] = -9'sd0;
	qsin_lut[105] = -9'sd150;
	icos_lut[105] =  9'sd30;
	qsin_lut[106] = -9'sd141;
	icos_lut[106] =  9'sd59;
	qsin_lut[107] = -9'sd127;
	icos_lut[107] =  9'sd85;
	qsin_lut[108] = -9'sd108;
	icos_lut[108] =  9'sd108;
	qsin_lut[109] = -9'sd85;
	icos_lut[109] =  9'sd127;
	qsin_lut[110] = -9'sd59;
	icos_lut[110] =  9'sd141;
	qsin_lut[111] = -9'sd30;
	icos_lut[111] =  9'sd150;
	qsin_lut[112] = -9'sd0;
	icos_lut[112] =  9'sd153;
	qsin_lut[113] =  9'sd30;
	icos_lut[113] =  9'sd150;
	qsin_lut[114] =  9'sd59;
	icos_lut[114] =  9'sd141;
	qsin_lut[115] =  9'sd85;
	icos_lut[115] =  9'sd127;
	qsin_lut[116] =  9'sd108;
	icos_lut[116] =  9'sd108;
	qsin_lut[117] =  9'sd127;
	icos_lut[117] =  9'sd85;
	qsin_lut[118] =  9'sd141;
	icos_lut[118] =  9'sd59;
	qsin_lut[119] =  9'sd150;
	icos_lut[119] =  9'sd30;
	qsin_lut[120] =  9'sd153;
	icos_lut[120] =  9'sd0;
	qsin_lut[121] =  9'sd150;
	icos_lut[121] = -9'sd30;
	qsin_lut[122] =  9'sd141;
	icos_lut[122] = -9'sd59;
	qsin_lut[123] =  9'sd127;
	icos_lut[123] = -9'sd85;
	qsin_lut[124] =  9'sd108;
	icos_lut[124] = -9'sd108;
	qsin_lut[125] =  9'sd85;
	icos_lut[125] = -9'sd127;
	qsin_lut[126] =  9'sd59;
	icos_lut[126] = -9'sd141;
	qsin_lut[127] =  9'sd30;
	icos_lut[127] = -9'sd150;
	qsin_lut[128] =  9'sd0;
	icos_lut[128] = -9'sd119;
	qsin_lut[129] = -9'sd23;
	icos_lut[129] = -9'sd117;
	qsin_lut[130] = -9'sd46;
	icos_lut[130] = -9'sd110;
	qsin_lut[131] = -9'sd66;
	icos_lut[131] = -9'sd99;
	qsin_lut[132] = -9'sd84;
	icos_lut[132] = -9'sd84;
	qsin_lut[133] = -9'sd99;
	icos_lut[133] = -9'sd66;
	qsin_lut[134] = -9'sd110;
	icos_lut[134] = -9'sd46;
	qsin_lut[135] = -9'sd117;
	icos_lut[135] = -9'sd23;
	qsin_lut[136] = -9'sd119;
	icos_lut[136] = -9'sd0;
	qsin_lut[137] = -9'sd117;
	icos_lut[137] =  9'sd23;
	qsin_lut[138] = -9'sd110;
	icos_lut[138] =  9'sd46;
	qsin_lut[139] = -9'sd99;
	icos_lut[139] =  9'sd66;
	qsin_lut[140] = -9'sd84;
	icos_lut[140] =  9'sd84;
	qsin_lut[141] = -9'sd66;
	icos_lut[141] =  9'sd99;
	qsin_lut[142] = -9'sd46;
	icos_lut[142] =  9'sd110;
	qsin_lut[143] = -9'sd23;
	icos_lut[143] =  9'sd117;
	qsin_lut[144] = -9'sd0;
	icos_lut[144] =  9'sd119;
	qsin_lut[145] =  9'sd23;
	icos_lut[145] =  9'sd117;
	qsin_lut[146] =  9'sd46;
	icos_lut[146] =  9'sd110;
	qsin_lut[147] =  9'sd66;
	icos_lut[147] =  9'sd99;
	qsin_lut[148] =  9'sd84;
	icos_lut[148] =  9'sd84;
	qsin_lut[149] =  9'sd99;
	icos_lut[149] =  9'sd66;
	qsin_lut[150] =  9'sd110;
	icos_lut[150] =  9'sd46;
	qsin_lut[151] =  9'sd117;
	icos_lut[151] =  9'sd23;
	qsin_lut[152] =  9'sd119;
	icos_lut[152] =  9'sd0;
	qsin_lut[153] =  9'sd117;
	icos_lut[153] = -9'sd23;
	qsin_lut[154] =  9'sd110;
	icos_lut[154] = -9'sd46;
	qsin_lut[155] =  9'sd99;
	icos_lut[155] = -9'sd66;
	qsin_lut[156] =  9'sd84;
	icos_lut[156] = -9'sd84;
	qsin_lut[157] =  9'sd66;
	icos_lut[157] = -9'sd99;
	qsin_lut[158] =  9'sd46;
	icos_lut[158] = -9'sd110;
	qsin_lut[159] =  9'sd23;
	icos_lut[159] = -9'sd117;
	qsin_lut[160] =  9'sd0;
	icos_lut[160] = -9'sd85;
	qsin_lut[161] = -9'sd17;
	icos_lut[161] = -9'sd83;
	qsin_lut[162] = -9'sd33;
	icos_lut[162] = -9'sd79;
	qsin_lut[163] = -9'sd47;
	icos_lut[163] = -9'sd71;
	qsin_lut[164] = -9'sd60;
	icos_lut[164] = -9'sd60;
	qsin_lut[165] = -9'sd71;
	icos_lut[165] = -9'sd47;
	qsin_lut[166] = -9'sd79;
	icos_lut[166] = -9'sd33;
	qsin_lut[167] = -9'sd83;
	icos_lut[167] = -9'sd17;
	qsin_lut[168] = -9'sd85;
	icos_lut[168] = -9'sd0;
	qsin_lut[169] = -9'sd83;
	icos_lut[169] =  9'sd17;
	qsin_lut[170] = -9'sd79;
	icos_lut[170] =  9'sd33;
	qsin_lut[171] = -9'sd71;
	icos_lut[171] =  9'sd47;
	qsin_lut[172] = -9'sd60;
	icos_lut[172] =  9'sd60;
	qsin_lut[173] = -9'sd47;
	icos_lut[173] =  9'sd71;
	qsin_lut[174] = -9'sd33;
	icos_lut[174] =  9'sd79;
	qsin_lut[175] = -9'sd17;
	icos_lut[175] =  9'sd83;
	qsin_lut[176] = -9'sd0;
	icos_lut[176] =  9'sd85;
	qsin_lut[177] =  9'sd17;
	icos_lut[177] =  9'sd83;
	qsin_lut[178] =  9'sd33;
	icos_lut[178] =  9'sd79;
	qsin_lut[179] =  9'sd47;
	icos_lut[179] =  9'sd71;
	qsin_lut[180] =  9'sd60;
	icos_lut[180] =  9'sd60;
	qsin_lut[181] =  9'sd71;
	icos_lut[181] =  9'sd47;
	qsin_lut[182] =  9'sd79;
	icos_lut[182] =  9'sd33;
	qsin_lut[183] =  9'sd83;
	icos_lut[183] =  9'sd17;
	qsin_lut[184] =  9'sd85;
	icos_lut[184] =  9'sd0;
	qsin_lut[185] =  9'sd83;
	icos_lut[185] = -9'sd17;
	qsin_lut[186] =  9'sd79;
	icos_lut[186] = -9'sd33;
	qsin_lut[187] =  9'sd71;
	icos_lut[187] = -9'sd47;
	qsin_lut[188] =  9'sd60;
	icos_lut[188] = -9'sd60;
	qsin_lut[189] =  9'sd47;
	icos_lut[189] = -9'sd71;
	qsin_lut[190] =  9'sd33;
	icos_lut[190] = -9'sd79;
	qsin_lut[191] =  9'sd17;
	icos_lut[191] = -9'sd83;
	qsin_lut[192] =  9'sd0;
	icos_lut[192] = -9'sd51;
	qsin_lut[193] = -9'sd10;
	icos_lut[193] = -9'sd50;
	qsin_lut[194] = -9'sd20;
	icos_lut[194] = -9'sd47;
	qsin_lut[195] = -9'sd28;
	icos_lut[195] = -9'sd42;
	qsin_lut[196] = -9'sd36;
	icos_lut[196] = -9'sd36;
	qsin_lut[197] = -9'sd42;
	icos_lut[197] = -9'sd28;
	qsin_lut[198] = -9'sd47;
	icos_lut[198] = -9'sd20;
	qsin_lut[199] = -9'sd50;
	icos_lut[199] = -9'sd10;
	qsin_lut[200] = -9'sd51;
	icos_lut[200] = -9'sd0;
	qsin_lut[201] = -9'sd50;
	icos_lut[201] =  9'sd10;
	qsin_lut[202] = -9'sd47;
	icos_lut[202] =  9'sd20;
	qsin_lut[203] = -9'sd42;
	icos_lut[203] =  9'sd28;
	qsin_lut[204] = -9'sd36;
	icos_lut[204] =  9'sd36;
	qsin_lut[205] = -9'sd28;
	icos_lut[205] =  9'sd42;
	qsin_lut[206] = -9'sd20;
	icos_lut[206] =  9'sd47;
	qsin_lut[207] = -9'sd10;
	icos_lut[207] =  9'sd50;
	qsin_lut[208] = -9'sd0;
	icos_lut[208] =  9'sd51;
	qsin_lut[209] =  9'sd10;
	icos_lut[209] =  9'sd50;
	qsin_lut[210] =  9'sd20;
	icos_lut[210] =  9'sd47;
	qsin_lut[211] =  9'sd28;
	icos_lut[211] =  9'sd42;
	qsin_lut[212] =  9'sd36;
	icos_lut[212] =  9'sd36;
	qsin_lut[213] =  9'sd42;
	icos_lut[213] =  9'sd28;
	qsin_lut[214] =  9'sd47;
	icos_lut[214] =  9'sd20;
	qsin_lut[215] =  9'sd50;
	icos_lut[215] =  9'sd10;
	qsin_lut[216] =  9'sd51;
	icos_lut[216] =  9'sd0;
	qsin_lut[217] =  9'sd50;
	icos_lut[217] = -9'sd10;
	qsin_lut[218] =  9'sd47;
	icos_lut[218] = -9'sd20;
	qsin_lut[219] =  9'sd42;
	icos_lut[219] = -9'sd28;
	qsin_lut[220] =  9'sd36;
	icos_lut[220] = -9'sd36;
	qsin_lut[221] =  9'sd28;
	icos_lut[221] = -9'sd42;
	qsin_lut[222] =  9'sd20;
	icos_lut[222] = -9'sd47;
	qsin_lut[223] =  9'sd10;
	icos_lut[223] = -9'sd50;
	qsin_lut[224] =  9'sd0;
	icos_lut[224] = -9'sd17;
	qsin_lut[225] = -9'sd3;
	icos_lut[225] = -9'sd17;
	qsin_lut[226] = -9'sd7;
	icos_lut[226] = -9'sd16;
	qsin_lut[227] = -9'sd9;
	icos_lut[227] = -9'sd14;
	qsin_lut[228] = -9'sd12;
	icos_lut[228] = -9'sd12;
	qsin_lut[229] = -9'sd14;
	icos_lut[229] = -9'sd9;
	qsin_lut[230] = -9'sd16;
	icos_lut[230] = -9'sd7;
	qsin_lut[231] = -9'sd17;
	icos_lut[231] = -9'sd3;
	qsin_lut[232] = -9'sd17;
	icos_lut[232] = -9'sd0;
	qsin_lut[233] = -9'sd17;
	icos_lut[233] =  9'sd3;
	qsin_lut[234] = -9'sd16;
	icos_lut[234] =  9'sd7;
	qsin_lut[235] = -9'sd14;
	icos_lut[235] =  9'sd9;
	qsin_lut[236] = -9'sd12;
	icos_lut[236] =  9'sd12;
	qsin_lut[237] = -9'sd9;
	icos_lut[237] =  9'sd14;
	qsin_lut[238] = -9'sd7;
	icos_lut[238] =  9'sd16;
	qsin_lut[239] = -9'sd3;
	icos_lut[239] =  9'sd17;
	qsin_lut[240] = -9'sd0;
	icos_lut[240] =  9'sd17;
	qsin_lut[241] =  9'sd3;
	icos_lut[241] =  9'sd17;
	qsin_lut[242] =  9'sd7;
	icos_lut[242] =  9'sd16;
	qsin_lut[243] =  9'sd9;
	icos_lut[243] =  9'sd14;
	qsin_lut[244] =  9'sd12;
	icos_lut[244] =  9'sd12;
	qsin_lut[245] =  9'sd14;
	icos_lut[245] =  9'sd9;
	qsin_lut[246] =  9'sd16;
	icos_lut[246] =  9'sd7;
	qsin_lut[247] =  9'sd17;
	icos_lut[247] =  9'sd3;
	qsin_lut[248] =  9'sd17;
	icos_lut[248] =  9'sd0;
	qsin_lut[249] =  9'sd17;
	icos_lut[249] = -9'sd3;
	qsin_lut[250] =  9'sd16;
	icos_lut[250] = -9'sd7;
	qsin_lut[251] =  9'sd14;
	icos_lut[251] = -9'sd9;
	qsin_lut[252] =  9'sd12;
	icos_lut[252] = -9'sd12;
	qsin_lut[253] =  9'sd9;
	icos_lut[253] = -9'sd14;
	qsin_lut[254] =  9'sd7;
	icos_lut[254] = -9'sd16;
	qsin_lut[255] =  9'sd3;
	icos_lut[255] = -9'sd17;
	qsin_lut[256] =  9'sd0;
	icos_lut[256] =  9'sd17;
	qsin_lut[257] =  9'sd3;
	icos_lut[257] =  9'sd17;
	qsin_lut[258] =  9'sd7;
	icos_lut[258] =  9'sd16;
	qsin_lut[259] =  9'sd9;
	icos_lut[259] =  9'sd14;
	qsin_lut[260] =  9'sd12;
	icos_lut[260] =  9'sd12;
	qsin_lut[261] =  9'sd14;
	icos_lut[261] =  9'sd9;
	qsin_lut[262] =  9'sd16;
	icos_lut[262] =  9'sd7;
	qsin_lut[263] =  9'sd17;
	icos_lut[263] =  9'sd3;
	qsin_lut[264] =  9'sd17;
	icos_lut[264] =  9'sd0;
	qsin_lut[265] =  9'sd17;
	icos_lut[265] = -9'sd3;
	qsin_lut[266] =  9'sd16;
	icos_lut[266] = -9'sd7;
	qsin_lut[267] =  9'sd14;
	icos_lut[267] = -9'sd9;
	qsin_lut[268] =  9'sd12;
	icos_lut[268] = -9'sd12;
	qsin_lut[269] =  9'sd9;
	icos_lut[269] = -9'sd14;
	qsin_lut[270] =  9'sd7;
	icos_lut[270] = -9'sd16;
	qsin_lut[271] =  9'sd3;
	icos_lut[271] = -9'sd17;
	qsin_lut[272] =  9'sd0;
	icos_lut[272] = -9'sd17;
	qsin_lut[273] = -9'sd3;
	icos_lut[273] = -9'sd17;
	qsin_lut[274] = -9'sd7;
	icos_lut[274] = -9'sd16;
	qsin_lut[275] = -9'sd9;
	icos_lut[275] = -9'sd14;
	qsin_lut[276] = -9'sd12;
	icos_lut[276] = -9'sd12;
	qsin_lut[277] = -9'sd14;
	icos_lut[277] = -9'sd9;
	qsin_lut[278] = -9'sd16;
	icos_lut[278] = -9'sd7;
	qsin_lut[279] = -9'sd17;
	icos_lut[279] = -9'sd3;
	qsin_lut[280] = -9'sd17;
	icos_lut[280] = -9'sd0;
	qsin_lut[281] = -9'sd17;
	icos_lut[281] =  9'sd3;
	qsin_lut[282] = -9'sd16;
	icos_lut[282] =  9'sd7;
	qsin_lut[283] = -9'sd14;
	icos_lut[283] =  9'sd9;
	qsin_lut[284] = -9'sd12;
	icos_lut[284] =  9'sd12;
	qsin_lut[285] = -9'sd9;
	icos_lut[285] =  9'sd14;
	qsin_lut[286] = -9'sd7;
	icos_lut[286] =  9'sd16;
	qsin_lut[287] = -9'sd3;
	icos_lut[287] =  9'sd17;
	qsin_lut[288] =  9'sd0;
	icos_lut[288] =  9'sd51;
	qsin_lut[289] =  9'sd10;
	icos_lut[289] =  9'sd50;
	qsin_lut[290] =  9'sd20;
	icos_lut[290] =  9'sd47;
	qsin_lut[291] =  9'sd28;
	icos_lut[291] =  9'sd42;
	qsin_lut[292] =  9'sd36;
	icos_lut[292] =  9'sd36;
	qsin_lut[293] =  9'sd42;
	icos_lut[293] =  9'sd28;
	qsin_lut[294] =  9'sd47;
	icos_lut[294] =  9'sd20;
	qsin_lut[295] =  9'sd50;
	icos_lut[295] =  9'sd10;
	qsin_lut[296] =  9'sd51;
	icos_lut[296] =  9'sd0;
	qsin_lut[297] =  9'sd50;
	icos_lut[297] = -9'sd10;
	qsin_lut[298] =  9'sd47;
	icos_lut[298] = -9'sd20;
	qsin_lut[299] =  9'sd42;
	icos_lut[299] = -9'sd28;
	qsin_lut[300] =  9'sd36;
	icos_lut[300] = -9'sd36;
	qsin_lut[301] =  9'sd28;
	icos_lut[301] = -9'sd42;
	qsin_lut[302] =  9'sd20;
	icos_lut[302] = -9'sd47;
	qsin_lut[303] =  9'sd10;
	icos_lut[303] = -9'sd50;
	qsin_lut[304] =  9'sd0;
	icos_lut[304] = -9'sd51;
	qsin_lut[305] = -9'sd10;
	icos_lut[305] = -9'sd50;
	qsin_lut[306] = -9'sd20;
	icos_lut[306] = -9'sd47;
	qsin_lut[307] = -9'sd28;
	icos_lut[307] = -9'sd42;
	qsin_lut[308] = -9'sd36;
	icos_lut[308] = -9'sd36;
	qsin_lut[309] = -9'sd42;
	icos_lut[309] = -9'sd28;
	qsin_lut[310] = -9'sd47;
	icos_lut[310] = -9'sd20;
	qsin_lut[311] = -9'sd50;
	icos_lut[311] = -9'sd10;
	qsin_lut[312] = -9'sd51;
	icos_lut[312] = -9'sd0;
	qsin_lut[313] = -9'sd50;
	icos_lut[313] =  9'sd10;
	qsin_lut[314] = -9'sd47;
	icos_lut[314] =  9'sd20;
	qsin_lut[315] = -9'sd42;
	icos_lut[315] =  9'sd28;
	qsin_lut[316] = -9'sd36;
	icos_lut[316] =  9'sd36;
	qsin_lut[317] = -9'sd28;
	icos_lut[317] =  9'sd42;
	qsin_lut[318] = -9'sd20;
	icos_lut[318] =  9'sd47;
	qsin_lut[319] = -9'sd10;
	icos_lut[319] =  9'sd50;
	qsin_lut[320] =  9'sd0;
	icos_lut[320] =  9'sd85;
	qsin_lut[321] =  9'sd17;
	icos_lut[321] =  9'sd83;
	qsin_lut[322] =  9'sd33;
	icos_lut[322] =  9'sd79;
	qsin_lut[323] =  9'sd47;
	icos_lut[323] =  9'sd71;
	qsin_lut[324] =  9'sd60;
	icos_lut[324] =  9'sd60;
	qsin_lut[325] =  9'sd71;
	icos_lut[325] =  9'sd47;
	qsin_lut[326] =  9'sd79;
	icos_lut[326] =  9'sd33;
	qsin_lut[327] =  9'sd83;
	icos_lut[327] =  9'sd17;
	qsin_lut[328] =  9'sd85;
	icos_lut[328] =  9'sd0;
	qsin_lut[329] =  9'sd83;
	icos_lut[329] = -9'sd17;
	qsin_lut[330] =  9'sd79;
	icos_lut[330] = -9'sd33;
	qsin_lut[331] =  9'sd71;
	icos_lut[331] = -9'sd47;
	qsin_lut[332] =  9'sd60;
	icos_lut[332] = -9'sd60;
	qsin_lut[333] =  9'sd47;
	icos_lut[333] = -9'sd71;
	qsin_lut[334] =  9'sd33;
	icos_lut[334] = -9'sd79;
	qsin_lut[335] =  9'sd17;
	icos_lut[335] = -9'sd83;
	qsin_lut[336] =  9'sd0;
	icos_lut[336] = -9'sd85;
	qsin_lut[337] = -9'sd17;
	icos_lut[337] = -9'sd83;
	qsin_lut[338] = -9'sd33;
	icos_lut[338] = -9'sd79;
	qsin_lut[339] = -9'sd47;
	icos_lut[339] = -9'sd71;
	qsin_lut[340] = -9'sd60;
	icos_lut[340] = -9'sd60;
	qsin_lut[341] = -9'sd71;
	icos_lut[341] = -9'sd47;
	qsin_lut[342] = -9'sd79;
	icos_lut[342] = -9'sd33;
	qsin_lut[343] = -9'sd83;
	icos_lut[343] = -9'sd17;
	qsin_lut[344] = -9'sd85;
	icos_lut[344] = -9'sd0;
	qsin_lut[345] = -9'sd83;
	icos_lut[345] =  9'sd17;
	qsin_lut[346] = -9'sd79;
	icos_lut[346] =  9'sd33;
	qsin_lut[347] = -9'sd71;
	icos_lut[347] =  9'sd47;
	qsin_lut[348] = -9'sd60;
	icos_lut[348] =  9'sd60;
	qsin_lut[349] = -9'sd47;
	icos_lut[349] =  9'sd71;
	qsin_lut[350] = -9'sd33;
	icos_lut[350] =  9'sd79;
	qsin_lut[351] = -9'sd17;
	icos_lut[351] =  9'sd83;
	qsin_lut[352] =  9'sd0;
	icos_lut[352] =  9'sd119;
	qsin_lut[353] =  9'sd23;
	icos_lut[353] =  9'sd117;
	qsin_lut[354] =  9'sd46;
	icos_lut[354] =  9'sd110;
	qsin_lut[355] =  9'sd66;
	icos_lut[355] =  9'sd99;
	qsin_lut[356] =  9'sd84;
	icos_lut[356] =  9'sd84;
	qsin_lut[357] =  9'sd99;
	icos_lut[357] =  9'sd66;
	qsin_lut[358] =  9'sd110;
	icos_lut[358] =  9'sd46;
	qsin_lut[359] =  9'sd117;
	icos_lut[359] =  9'sd23;
	qsin_lut[360] =  9'sd119;
	icos_lut[360] =  9'sd0;
	qsin_lut[361] =  9'sd117;
	icos_lut[361] = -9'sd23;
	qsin_lut[362] =  9'sd110;
	icos_lut[362] = -9'sd46;
	qsin_lut[363] =  9'sd99;
	icos_lut[363] = -9'sd66;
	qsin_lut[364] =  9'sd84;
	icos_lut[364] = -9'sd84;
	qsin_lut[365] =  9'sd66;
	icos_lut[365] = -9'sd99;
	qsin_lut[366] =  9'sd46;
	icos_lut[366] = -9'sd110;
	qsin_lut[367] =  9'sd23;
	icos_lut[367] = -9'sd117;
	qsin_lut[368] =  9'sd0;
	icos_lut[368] = -9'sd119;
	qsin_lut[369] = -9'sd23;
	icos_lut[369] = -9'sd117;
	qsin_lut[370] = -9'sd46;
	icos_lut[370] = -9'sd110;
	qsin_lut[371] = -9'sd66;
	icos_lut[371] = -9'sd99;
	qsin_lut[372] = -9'sd84;
	icos_lut[372] = -9'sd84;
	qsin_lut[373] = -9'sd99;
	icos_lut[373] = -9'sd66;
	qsin_lut[374] = -9'sd110;
	icos_lut[374] = -9'sd46;
	qsin_lut[375] = -9'sd117;
	icos_lut[375] = -9'sd23;
	qsin_lut[376] = -9'sd119;
	icos_lut[376] = -9'sd0;
	qsin_lut[377] = -9'sd117;
	icos_lut[377] =  9'sd23;
	qsin_lut[378] = -9'sd110;
	icos_lut[378] =  9'sd46;
	qsin_lut[379] = -9'sd99;
	icos_lut[379] =  9'sd66;
	qsin_lut[380] = -9'sd84;
	icos_lut[380] =  9'sd84;
	qsin_lut[381] = -9'sd66;
	icos_lut[381] =  9'sd99;
	qsin_lut[382] = -9'sd46;
	icos_lut[382] =  9'sd110;
	qsin_lut[383] = -9'sd23;
	icos_lut[383] =  9'sd117;
	qsin_lut[384] =  9'sd0;
	icos_lut[384] =  9'sd153;
	qsin_lut[385] =  9'sd30;
	icos_lut[385] =  9'sd150;
	qsin_lut[386] =  9'sd59;
	icos_lut[386] =  9'sd141;
	qsin_lut[387] =  9'sd85;
	icos_lut[387] =  9'sd127;
	qsin_lut[388] =  9'sd108;
	icos_lut[388] =  9'sd108;
	qsin_lut[389] =  9'sd127;
	icos_lut[389] =  9'sd85;
	qsin_lut[390] =  9'sd141;
	icos_lut[390] =  9'sd59;
	qsin_lut[391] =  9'sd150;
	icos_lut[391] =  9'sd30;
	qsin_lut[392] =  9'sd153;
	icos_lut[392] =  9'sd0;
	qsin_lut[393] =  9'sd150;
	icos_lut[393] = -9'sd30;
	qsin_lut[394] =  9'sd141;
	icos_lut[394] = -9'sd59;
	qsin_lut[395] =  9'sd127;
	icos_lut[395] = -9'sd85;
	qsin_lut[396] =  9'sd108;
	icos_lut[396] = -9'sd108;
	qsin_lut[397] =  9'sd85;
	icos_lut[397] = -9'sd127;
	qsin_lut[398] =  9'sd59;
	icos_lut[398] = -9'sd141;
	qsin_lut[399] =  9'sd30;
	icos_lut[399] = -9'sd150;
	qsin_lut[400] =  9'sd0;
	icos_lut[400] = -9'sd153;
	qsin_lut[401] = -9'sd30;
	icos_lut[401] = -9'sd150;
	qsin_lut[402] = -9'sd59;
	icos_lut[402] = -9'sd141;
	qsin_lut[403] = -9'sd85;
	icos_lut[403] = -9'sd127;
	qsin_lut[404] = -9'sd108;
	icos_lut[404] = -9'sd108;
	qsin_lut[405] = -9'sd127;
	icos_lut[405] = -9'sd85;
	qsin_lut[406] = -9'sd141;
	icos_lut[406] = -9'sd59;
	qsin_lut[407] = -9'sd150;
	icos_lut[407] = -9'sd30;
	qsin_lut[408] = -9'sd153;
	icos_lut[408] = -9'sd0;
	qsin_lut[409] = -9'sd150;
	icos_lut[409] =  9'sd30;
	qsin_lut[410] = -9'sd141;
	icos_lut[410] =  9'sd59;
	qsin_lut[411] = -9'sd127;
	icos_lut[411] =  9'sd85;
	qsin_lut[412] = -9'sd108;
	icos_lut[412] =  9'sd108;
	qsin_lut[413] = -9'sd85;
	icos_lut[413] =  9'sd127;
	qsin_lut[414] = -9'sd59;
	icos_lut[414] =  9'sd141;
	qsin_lut[415] = -9'sd30;
	icos_lut[415] =  9'sd150;
	qsin_lut[416] =  9'sd0;
	icos_lut[416] =  9'sd187;
	qsin_lut[417] =  9'sd36;
	icos_lut[417] =  9'sd183;
	qsin_lut[418] =  9'sd72;
	icos_lut[418] =  9'sd173;
	qsin_lut[419] =  9'sd104;
	icos_lut[419] =  9'sd155;
	qsin_lut[420] =  9'sd132;
	icos_lut[420] =  9'sd132;
	qsin_lut[421] =  9'sd155;
	icos_lut[421] =  9'sd104;
	qsin_lut[422] =  9'sd173;
	icos_lut[422] =  9'sd72;
	qsin_lut[423] =  9'sd183;
	icos_lut[423] =  9'sd36;
	qsin_lut[424] =  9'sd187;
	icos_lut[424] =  9'sd0;
	qsin_lut[425] =  9'sd183;
	icos_lut[425] = -9'sd36;
	qsin_lut[426] =  9'sd173;
	icos_lut[426] = -9'sd72;
	qsin_lut[427] =  9'sd155;
	icos_lut[427] = -9'sd104;
	qsin_lut[428] =  9'sd132;
	icos_lut[428] = -9'sd132;
	qsin_lut[429] =  9'sd104;
	icos_lut[429] = -9'sd155;
	qsin_lut[430] =  9'sd72;
	icos_lut[430] = -9'sd173;
	qsin_lut[431] =  9'sd36;
	icos_lut[431] = -9'sd183;
	qsin_lut[432] =  9'sd0;
	icos_lut[432] = -9'sd187;
	qsin_lut[433] = -9'sd36;
	icos_lut[433] = -9'sd183;
	qsin_lut[434] = -9'sd72;
	icos_lut[434] = -9'sd173;
	qsin_lut[435] = -9'sd104;
	icos_lut[435] = -9'sd155;
	qsin_lut[436] = -9'sd132;
	icos_lut[436] = -9'sd132;
	qsin_lut[437] = -9'sd155;
	icos_lut[437] = -9'sd104;
	qsin_lut[438] = -9'sd173;
	icos_lut[438] = -9'sd72;
	qsin_lut[439] = -9'sd183;
	icos_lut[439] = -9'sd36;
	qsin_lut[440] = -9'sd187;
	icos_lut[440] = -9'sd0;
	qsin_lut[441] = -9'sd183;
	icos_lut[441] =  9'sd36;
	qsin_lut[442] = -9'sd173;
	icos_lut[442] =  9'sd72;
	qsin_lut[443] = -9'sd155;
	icos_lut[443] =  9'sd104;
	qsin_lut[444] = -9'sd132;
	icos_lut[444] =  9'sd132;
	qsin_lut[445] = -9'sd104;
	icos_lut[445] =  9'sd155;
	qsin_lut[446] = -9'sd72;
	icos_lut[446] =  9'sd173;
	qsin_lut[447] = -9'sd36;
	icos_lut[447] =  9'sd183;
	qsin_lut[448] =  9'sd0;
	icos_lut[448] =  9'sd221;
	qsin_lut[449] =  9'sd43;
	icos_lut[449] =  9'sd217;
	qsin_lut[450] =  9'sd85;
	icos_lut[450] =  9'sd204;
	qsin_lut[451] =  9'sd123;
	icos_lut[451] =  9'sd184;
	qsin_lut[452] =  9'sd156;
	icos_lut[452] =  9'sd156;
	qsin_lut[453] =  9'sd184;
	icos_lut[453] =  9'sd123;
	qsin_lut[454] =  9'sd204;
	icos_lut[454] =  9'sd85;
	qsin_lut[455] =  9'sd217;
	icos_lut[455] =  9'sd43;
	qsin_lut[456] =  9'sd221;
	icos_lut[456] =  9'sd0;
	qsin_lut[457] =  9'sd217;
	icos_lut[457] = -9'sd43;
	qsin_lut[458] =  9'sd204;
	icos_lut[458] = -9'sd85;
	qsin_lut[459] =  9'sd184;
	icos_lut[459] = -9'sd123;
	qsin_lut[460] =  9'sd156;
	icos_lut[460] = -9'sd156;
	qsin_lut[461] =  9'sd123;
	icos_lut[461] = -9'sd184;
	qsin_lut[462] =  9'sd85;
	icos_lut[462] = -9'sd204;
	qsin_lut[463] =  9'sd43;
	icos_lut[463] = -9'sd217;
	qsin_lut[464] =  9'sd0;
	icos_lut[464] = -9'sd221;
	qsin_lut[465] = -9'sd43;
	icos_lut[465] = -9'sd217;
	qsin_lut[466] = -9'sd85;
	icos_lut[466] = -9'sd204;
	qsin_lut[467] = -9'sd123;
	icos_lut[467] = -9'sd184;
	qsin_lut[468] = -9'sd156;
	icos_lut[468] = -9'sd156;
	qsin_lut[469] = -9'sd184;
	icos_lut[469] = -9'sd123;
	qsin_lut[470] = -9'sd204;
	icos_lut[470] = -9'sd85;
	qsin_lut[471] = -9'sd217;
	icos_lut[471] = -9'sd43;
	qsin_lut[472] = -9'sd221;
	icos_lut[472] = -9'sd0;
	qsin_lut[473] = -9'sd217;
	icos_lut[473] =  9'sd43;
	qsin_lut[474] = -9'sd204;
	icos_lut[474] =  9'sd85;
	qsin_lut[475] = -9'sd184;
	icos_lut[475] =  9'sd123;
	qsin_lut[476] = -9'sd156;
	icos_lut[476] =  9'sd156;
	qsin_lut[477] = -9'sd123;
	icos_lut[477] =  9'sd184;
	qsin_lut[478] = -9'sd85;
	icos_lut[478] =  9'sd204;
	qsin_lut[479] = -9'sd43;
	icos_lut[479] =  9'sd217;
	qsin_lut[480] =  9'sd0;
	icos_lut[480] =  9'sd255;
	qsin_lut[481] =  9'sd50;
	icos_lut[481] =  9'sd250;
	qsin_lut[482] =  9'sd98;
	icos_lut[482] =  9'sd236;
	qsin_lut[483] =  9'sd142;
	icos_lut[483] =  9'sd212;
	qsin_lut[484] =  9'sd180;
	icos_lut[484] =  9'sd180;
	qsin_lut[485] =  9'sd212;
	icos_lut[485] =  9'sd142;
	qsin_lut[486] =  9'sd236;
	icos_lut[486] =  9'sd98;
	qsin_lut[487] =  9'sd250;
	icos_lut[487] =  9'sd50;
	qsin_lut[488] =  9'sd255;
	icos_lut[488] =  9'sd0;
	qsin_lut[489] =  9'sd250;
	icos_lut[489] = -9'sd50;
	qsin_lut[490] =  9'sd236;
	icos_lut[490] = -9'sd98;
	qsin_lut[491] =  9'sd212;
	icos_lut[491] = -9'sd142;
	qsin_lut[492] =  9'sd180;
	icos_lut[492] = -9'sd180;
	qsin_lut[493] =  9'sd142;
	icos_lut[493] = -9'sd212;
	qsin_lut[494] =  9'sd98;
	icos_lut[494] = -9'sd236;
	qsin_lut[495] =  9'sd50;
	icos_lut[495] = -9'sd250;
	qsin_lut[496] =  9'sd0;
	icos_lut[496] = -9'sd255;
	qsin_lut[497] = -9'sd50;
	icos_lut[497] = -9'sd250;
	qsin_lut[498] = -9'sd98;
	icos_lut[498] = -9'sd236;
	qsin_lut[499] = -9'sd142;
	icos_lut[499] = -9'sd212;
	qsin_lut[500] = -9'sd180;
	icos_lut[500] = -9'sd180;
	qsin_lut[501] = -9'sd212;
	icos_lut[501] = -9'sd142;
	qsin_lut[502] = -9'sd236;
	icos_lut[502] = -9'sd98;
	qsin_lut[503] = -9'sd250;
	icos_lut[503] = -9'sd50;
	qsin_lut[504] = -9'sd255;
	icos_lut[504] = -9'sd0;
	qsin_lut[505] = -9'sd250;
	icos_lut[505] =  9'sd50;
	qsin_lut[506] = -9'sd236;
	icos_lut[506] =  9'sd98;
	qsin_lut[507] = -9'sd212;
	icos_lut[507] =  9'sd142;
	qsin_lut[508] = -9'sd180;
	icos_lut[508] =  9'sd180;
	qsin_lut[509] = -9'sd142;
	icos_lut[509] =  9'sd212;
	qsin_lut[510] = -9'sd98;
	icos_lut[510] =  9'sd236;
	qsin_lut[511] = -9'sd50;
	icos_lut[511] =  9'sd250;
end

always @(t,i,q)
	begin
		icos_addr=(i<<5)+t;
		qsin_addr=(q<<5)+t;
	end

endmodule
